../../TRUE_DUAL_PORT_RAM/rtl/true_dual_port_ram.sv