../../WINDOW_SLIDE/rtl/window_slide_wrapper.sv