../../CALCULATORUNIT/rtl/AccelCoreL1.vhd