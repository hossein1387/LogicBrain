../../CALCULATORUNIT/rtl/LineBufferL1.vhd