../../LINE_BUFFER/rtl/line_buffer.sv