../../CALCULATORUNIT/rtl/CalculatorUnit.vhd