../../CALCULATORUNIT/rtl/LineBufferL2.vhd