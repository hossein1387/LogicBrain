../../CONTROLLER/rtl/controller.sv