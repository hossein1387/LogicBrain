../../WINDOW_SLIDE/rtl/window_slide.sv