logic[511:0]weight_l1[1023:0]={512'b11001101011101000000000100001100000000111100000000010001111100001100001100001100111111001100110000000111001100000000010011110100001111010100010101110101000100010001001101010111001100000101111100110101001100000000110000010101000101001100000101110011010000010100110000110101111100110100000001010001000001000111000100000101001100110001000100000000000001111100010000000100000001111111110001111101010111011111001111110111111111010101010100110011001100011111110111110000011101010111110000111101110001000011001111000001,512'b11000100110101110001010111001101010000000011001101010011010001010000011100001100110000110011000000001101000000110011010101001100110001010111000100011101011111011100011101111101000001010001000000000001000100110000000111000101011100000011110011000000010011000101000011000011000001000011010011000001111100000101010101110101110111010011000100001111010100110111110011000111001101001100010011110000001101011101110001010011011100110100010001000100011100111100010011000000010101011100110000000100001101110011010001000001,512'b11110111000000000111000000001100110011010001000100010000010000001100010011011101000011011100011100000111000000010100110011111101000101000000110111010000001111010111110000000101001111000011111101011100000011010100000101110000111101000100000000110011010101001100010101011100010011111100000000000100111111111100010001001101000000000100010000010000010001010000001111000011000100110100110001000100010011001100110111011111010011011100010011010111110001110011111111110011010111110011010011000011000000110100111100000000,512'b00011101110101000111111100010000110001000100110011010011110000110111000100110011110100011100000111000000111100011101010001010000000100001100010101011100111100110100010100111111000111010011110101011101110100001100000101110101010000110101110001010101110111111100110000001100001111111100001111110011000000010111110011011100011100110001110011000001000111110001111111110111011111010100010111010100110101010101010101110100001100000000110001110000010000000101111101000011000000000100010100000100000101000101111100000101,512'b01001100000001001100011111000001010111001111000000000000011111010011110111010100010001111101011101111101000111000001001100111101010000000111010111111101000100110001010101111100000000110100001101011100011101000100010000010101111101000011111111011101000011000100010100011111110000001111010000110011010100011111110000111111000000001100000101110011011111001111000001110100001111001101110111111100000100000011010000111101010011000111011101010100110011010001011101010101111111010011001111000011010101010111000000111101,512'b01010101000000111111000101111111111101011111011101110011010000000100001101110100010000011101011101010101000011000000110000010011010001001100000001011100110111011101110111111101011111000101111100010001000001000101010101001111010011001111110101010001000001110000110001110000111111010000010100001101000011000100000101011100010000000011110000111101110001000000110000001101000000110100111100011101011101000011110000001101010000001111110000110000010000110001000000010000010000010101111101000100010100000111010011011100,512'b11010101111111110000111101011100010100001101000001010001011101110111010000110001010001010111110011010011010000010001010000000111010100111101000100000000010000011111001101011101001111000000000100000100011101001101010100010011000101000101011100110011000011111111001111001101000101001111010001110001001101010001010000010000011100011100111101000101110100010001110100110101000000010100111111110101000111000101001111000111000001110001001100010111000001010100011100001101111111000100001100010000110100000000000001010000,512'b01011100011100010100111111000101000101111111010000000011111100110111010000001100110000010111110011111100000001110001001111000011001101000011010011011100111101111100110100011100000100010011001111011101111100111111000001000000011101000000000100000001001100010101000000000111010001110000010111110001010011000100000101110101001100110100011111001101000011111111000111000111111111110000000001000011110000011101001100001101110001111100011100010001110100110101110101010111001100010101000000001100000001000100111111111100,512'b00010100110100000101010000000000000100011101001101011100110101011111110000001100000000110001110000001111000101110100110100010000000101110100010111110111111101110111110111001100010000011101001111111101010100000011001101010111110001110101110011000111010000010001011100010011000000010001111111111111001111000100111101001101000011000000010111110011010000111100000100111100011100110000000111010011010000010111001100000001010111000000111111110000110100110100111101110101001101011101011100110000000111010111010001010100,512'b00010001110111010000111100010111000111000100001100000001010111110011111111000000000001111100000000010000010101011101000011010000000100011111001100010111010001000000000100111101000111000001001100111111110011111100001111000011111100010001001100010101111100001100000000000001010000001101011101110000010011011100000100010100001100010111000101011100010111000101001111000000010000001100010111011100001101000111010000000111000001011111000011010000010011000000010001001100010001111100000111010100110101011111010000000100,512'b11000011001111001100010001111111001111111101011101111100110011000011010011001111110000001101010011000101000000110001000111010000000100110001110011110101001100000000111101010100000011011111000100111101111111110111011100001101000101000011111100000000010000010100001111010000010100011100001111011111000001010001110001110000000111000101001111110111000011110011011100010111011101001101010100000000000000000111110101000001000100110000110001011100001100001101011101111101011101000111000100000000001100111101001100110100,512'b00011101000011001101000000011101000100111100110101010000110001000100010100010001001100110001000111011101010100000000000101111100111100011101010011011111110000000100011111000000110100111111110000110101000011110000001101010111110011000100110011000100111101000001001100010101010011010001111111111111011101010100110000000100011111110011010011000100111100010011000100110111001111010000011111010011001101010101011100001101110011001100010001001101000011111100110000000001110111110001000000110111000100010111111111010000,512'b11010111000101010100000101010111110101011111001111000000110000001100110111010001000111111100000100010001111111001100110100010101001111010100000011000011001101001101001101000100011111001100111111111101001100110011000001111100110111001111000101010101000000000101111111000000011100000000110000011101000111000101110111111111000011011100001100000000010100110001000101000111110011110000000001010000111101001111111100010101011100110000110101001100001100001111110100110111110111010100000000000001011100000000000101000100,512'b11110100111101010011111101000111010001111100010111111100010111011100110000110111000011110000111101000000011111000001010100111101000001000011001111011100000011110100010000111111001100000011010011010100110101110011000001010000110111000001000100011111110100000000011111001101001100000101001101000100010001111111001111001100000011010011000111111101111101000001001101001100111101011100000000110111000001010100110000011101000111000111110100110100000001000011110100011100000111110011000000110001110011110011011111000111,512'b11010100001101000101000011010101010111110011010111011101000100000001000100000100000001111111000111111101111111000000011111010101000101111100010000011111000100000001011100010000000111000001001100010000001100001101001111000101011111000001010000110111110101111100111101010001011101010000011100000101010101000101110111000000010000111101110111010000110011000111010001111101010111000011000011001100001111110111110000000011011111111101111100010000000011001100011100010111011101010011000011110011000000000111110111000000,512'b00000011110000000001000001111111010101010011010111000101011100110111000001111101111101010101010011001101110100011111110101000101110100011101110000111111001100011101111101001100001100010000000000111111011100000000010001010011010001001100001100011100110011111100001100000100000000010000110011001111111101001111110000000011110001000011010001111111010011110100010000111101110111000001110111000101110000000101010000110111110100000001000001001111111100000111011111110100000100000111111101000011110000110000000100000001,512'b00110100000000110100010100000101001111010101111101001101000100000000111100111101010001011101110111001100010000000100111101010011010111000101000100010100001101110111110100000001011101010001000101110100001100001111010000110101011101000001110100110111111100111100010000010011000101000101110000001100010111000101011100001100000100110100000000110111010101000111000101010111110100110011000100001111000000000000110100001111111111010111010011000000110100011100000100111111111101000000000000001100010011000011010100001111,512'b00010101010011000011001101000101000100010100000100001100110000001101001100110001110001000111001101000101110101011100110100010111110001110101010100011101010000010100010101111100010101001100000000000101011100110100110001001100011100010011110100110000010000001101010011000011010101000011000100000001000111010111000111111100000101000100000011000011110100111111010011110100110001000101011101001101000011111101111100110111010100001100110100010101000001001100010100001101000100011101010000111101110011001111001100000111,512'b11000001010100001101010001000000000011000111001111011111000100110011011111000011000000111100001100111100010000001101011100110001111100110100011101001101010101111100000011110000011111110100001100010100111111000011110000110100000001111100111111011100110011110111000001110011000000000101111101110000010001010100010101010000010001000111111100110000001100001100000001000101110100110100000000110101001100110111000111010011110100011101000111010100000100111101000101010111011101000001000100111101001101010100011101010000,512'b00001101010000000100110011010000000100110011111111010101110100110111110100000011010000010011011111011101010101010011111101001111001111110000000000000011111100000000010000010100010101110111011100001100111111010101000101000001001100010100110100001100000011111111000111001111000111010001001100111101111101001101010000000111110111000100000000010100000011011100110101000100010101111100010000110001000100010001110000000000111111110100000000110000010000010000000000110111110011010001110100011101010101001101001111010100,512'b01000011000001000100001100000000011111010001000011001111000100110011011111110000000011001111000101011111111111111100010011110001010101000100010000011101011100010000111111110101000111010000110101001100011100110001010011000011111111110100110001011100000100000000110011111111000100010101010111110001000100110100000100000111000011110011000101011111010100010111000000011100110101000100001100010100000011010101110011011101000111110001110000010111110011010111110011110011110011110001000001011100000011011111000011110100,512'b00000000001111000000011101000011000001010000011101111100110111010011011111111101111100010001001100110111110100000111010111010100001101111101010100001111011111110100110000010111010000110111000100011111000011000101001101000000010011110101001111010100010101010101000111000100000000000101001100000000110101011101110000110101000100001111110011000100001111111100010001000011011111000011110001110000011100110011000011110101011111000111110101001111010100010001111111000011000000001101000101000001000000000101110101010100,512'b01111100000011110111110111010000011111010101110100110001110111010111111100011111110001001100010100010100010011110000000101111101010000010101111111011111000011110100111101000100110101111111010011010000111101000011000011001100000111111101000100110100111100111100000100111111001111110001110000000100110011001100000011000001011101111101000000000101010101000011001100110101000111000111000101110101000011010100010111000000000101000000010111110001011111000001110111001111110001000100010100011111001100010100000000000000,512'b00001100011101010011000100000001001111110011111111000100010011010000000100000100010001111100000100000101011100000101111111000000010000011111110001010100000111000111000100110111110100000101110000001111011100000000111111011111011100001111011100010011000011000000001100010100000101111100110111010111000000110101110101110011111100000100110100010111011111110001001100011101111101111111010000000100010111010011000100001100000000001111000001000001010001010101110101111100010001110111000011111111010011110101011101011101,512'b11111100110101111100010011111101000011111111110101110000110011111101000000000101010111110111010011011101011100110101010011000011001111000011000000000101010101001111010000110111110000011100011100000011000101011100110100110100111100000001000000110000110100010001010100001111110111000111111111010101110100010001111100011101110111110000000000010001000000010111110000010100010111000011011100010111011101111101110100111100110100010011000000111100110001110001010111001100000100000100000101011100111111000100000011111100,512'b01000101001101000000000001110001000001111100110001000011111101110111001100010011110101000111111101010101011100010101110011001100110011010111001111001100001101110000111111110000000101110111111111010000000000111100010011000011110000111101110011001111010011010101110101110111001100110111000111110000110111111100010011010100010011001101000100001101000100000100000100110011010101000011010100010001011100000111110000110101010011001101000011001100111100011100010011000100011111110100000011001100110100011100110000010011,512'b11000011000011010101110011000111110100010011000000000100000100001100000001000101001111000011000011000011000100110011000011010111111100011111011100011101110011110100110011010111110000000011000001000101000100111111010100000101110111011111110100010101000111000000110100110011011100000101110100010111110111010100000011010101000000011100111101010001000100011100001101001100110000011101011101011101110100010011011100001101011100001111001101110000001100000101000011010111001100110011011101010001011100000111110100001101,512'b11000000110011000000110011001100000000010111001111111101110000001111110000010011110100000000001111010000010001001100001111011111111111000001010101010011111111000001000000011100111100000000110111011111010100001101111101010111001111011100011111011111010000010101110000111101010001110111011100000100000000001111010000000011010000001111000001011111010011110111000001110011000000001100111111010101010001010011010100000101011100011111000001000100110101000100011111111100001100110001011111110001110011110001010011110100,512'b11000000111111000101011111000111110001010001001111010000011100111100110011000111010000111101010001110001011101010001011100000001011111000100110001000101010011110101000001001100000001110001000111000101111100000011001100011111000011001111000011010011110111111100010101010000010000010000011101110011010101001111010100000011000111010001110100010101110011001100001111110001010111000101010011010001110101111111010100111100110100111101011101110111001101001101011101111111000000111111000011010011110011110000111100111101,512'b01001100110111010100110100000011000011110000000000111111011100011111000100010001110000111101000011111101010100010001010011111100110100000001110011010000001100000101110011110000110000000111001100110011010101010111110011011111010111111111011100110101110101110000001111010001111101010111110001111111110000111100110101001101010100000101110100110100000100010001000011001101000001001111010000110100010011000000010101010000110011001100110111011111000100001100000000000000000111111101110000110011011111010000011101000001,512'b01001111010001110001111111001100011100110000000100111100110100110101011100010011111100110100110000001111110000111101110011011111000000010100000001001111110001010000110011000100111100000111110000111111000011010000000001110100110100000000000000001100000011010100110111010000110000010100010100111100110111000111001101010001110000000100110100000011000000010000011101111101010100111111001100011100110100000000110100010100010001111101000101001111111100000001110000110001010111001101001100000101110001000001110100110111,512'b00011100010011000000000101110100000000000100110111010111000000110100010011010011110100110000001100001100110100000101110001110001000111010100010100011111000001011111000000010001110000000111011100010011110100000001000000001100111100110111000111010101010101000011010011111100000101010100110101111111001101010111001100011100001100010011000011000011001111001101110000000001000111000000010000111100111101011111011111010100001101010001110101001111000011000011000001001100111101110011000001110000010111000001010101110000,512'b01111111000001110000010111011101110100010000110101111111000100000011110100110000000000010100011100010111000011110101010000111111010000110100010100010100001100001100010100111100111100000101111100111101111111111101010000001100000101110011111111110000110101111101110101000001010001110001010101001101110100110100000100000111111101110000110000110101111101110001010000001100110101110000110101010100000001110011010101000001010101000100001101010100000011000100000101000011011111011100000100011101001111001100111111001111,512'b00110000001111000101010001001111010000010111110111000000110001011111010001111101001101010100010011110011110100001101010100111111010100000000000000110101000100001100000001110101110101000001001101010001010000010011001100110101011111111111000001000000010001001100110100001111011111001101110000010111110100111111011101010001011111110100010000110100110001000000000001110100001111010100010000001100011100110111010011010011111100111101010011110000000101001111110001001111011100110111110011110100010111000101110101110011,512'b11110111011100001100110001010011010011010001111100010101011100010100010101010001110000000100010001110000010111011111110100000111000111010001110011110111000111111100000011000100001111110111110001000011111100000000010000011111110000110100001100110011000001110001001101010011010100000100111111010011010011010011010100110100111100010101000111110000110100000000110111110111000011000111000100111100110011110001111100011101010001000011110100110001110001110101110000110001010011000101111101000101010111110100010100110011,512'b11110011010100011101001101110000111100010001110000000011110100000011110101001100111100001101001111110000011101010111010011111101110101001101011111010000110000111100110011110100000011010000010101010001011111000100011100110101010000110000000001001100000100000001000111110100011100010111010001111100010011001111011111011100011100000000000100110101000011010011011100011100010000111100000111110001110001000000010000010011001111010001000011010100111111111111110000011111000111011111010101000111111100010011110100110000,512'b01111101110000110000110000010001010000111101000001000000011111110011010000000000010101000001000111000100001100001100001100010111001111011101010111110011010011010001000011010011111101010001010000001111010100010000111101010001110001010011110011000000000100010011010000110011010100011100010011010000110000111111011101001111110111001100110111000101010100110001001100000011110000000011110101110000110100000000001100010011110001011100000111010100000101110000110101000011000000111101000011010001000101000100010111000000,512'b11010000000001001111110011011101011111010000001101110111110011010111001101010111110011000100011100000100000111111111110000010100000100011100010000010001011111010011000001110011110111011111000011000101010111010011011100000101000011000001000100011100010101010000000111110101010011000000111111111111000000110011110011001111010000011101001100000011000000111100111111001100010111110100000111000101000100010011011101011100010001011101001111110000010100010001010111010000010000000111000000011111110100110111001111010000,512'b00011111010101110101000100011111000111000001000001010011000001110100110111000101111100010100001100110011110001000100010001000100010011010000000011000100110001010111110000110011000101010000110001001100010011010000000100010100001100000011000101000000000101000000010001000100001101000000010011000011110111011101001100110000000101010001110000011101000100000000001100110111111111010111110111110111000000000001000011000101111111000111000011011111010000010011111100110000000101011111011100000111001101010000010001010100,512'b01010111010111111100010101010000110101000001000100011101001100110011000000010011000100001101000100011111110100110100000101000001110000110000010101001100011111010101001100111111110011000111110001110100000011001100110111110000011111001111010011010100110011010100110100001101000001010100111100000100000001110011111100000101110001111100000111110111010111111101010111000101110001000101110011110101001111000000010100011100011101001100110001000100111100010111111100110001010000010000111111010101010001010111010001010011,512'b00010001000100110000010011000111000101110111010100010101000011001101000101010000010101010001110001110100110101000101111101111100011100000000011111010001010100000001000000111100010001000011000011000011000001010011011101111100110101010011010000001100000100000011001101010101011101010111110111010000110000010100011100000101001111000111001101000101111101110100000011010101110111000011110111010011000001111100010101010111000000000000010100010101111100111100110100010000000101000000110000010001000101000001011111010000,512'b00000100011100111100011111111101010100110001010111001100001101010101110000110111111101000001001101011100000000010001111100110111010101000000110011000011011111000101011111010000011111110001000101000011010001000101110101001111111101000011110001010101000000111100011100001100111100110111000000110100010001001101110000111111001100001101110011010101000111000001010000010111000111011101011101001100111111011100110000110001011111111111110011001100110100010101000100001101001100110101110101010101010101011111000101001111,512'b11110101001100000101110001011111000101010001001111110011010100000011000001010111000001001101111101110000010101110100110111010101000101110001010001111111001111000000011101010000011101000001000100010101010100010011010100000101010011001100011100001100111101000111000100110011001111010111000000000011000111000100110000000001010100000101110000010100000101110000110101110001110011010000110101000011000111010011110000110001010001111100000101110100111111000100000001000100011101111100011111000000001100000111010011110100,512'b11001100110111000100110111011101010000110111000001010101110101000011110000010111000011000101000101000011001100110111110111001111000011001111011111001100010000110111111100110000111100000001111100000101000011111100000111110101110111000011001101000001000001000000010011110011001100010001000011110100110011110001000101111101010001110101010101000000011101110000010111011100010011000000000111110100000011000111010000110000000000001111010011110001110111011100010011000111000001000101110100110000001100110000000011110011,512'b00011101001100000100010001010001001101000111000000011101111100110011110100110100011100000111010100110011010101011101001101001101000001000011010011110001111101010000110011110011110101000001111101001101010111011111000111110111110000001100000100010000110000110100000100001111111100000001110011001100110100000101110111111111110001111100000100110000111101110100000011111100010011000100001100001111110011000011000101111111010001000011010100110000011111001100111111001101010000110100000101111100110011000000111111000001,512'b01001111110101001111000100110000011101110111010111000111110000000001010000010001110100010100010000010001010111010101010000000001111101010011010000110100010000000101110001010100000000010101010011010000001100000101111111000100001100000001000100111111011101111101010001110011001100011111000011111101110100110101110101110000011111111100001111010001010000001100000011010000110100111101011100111101001101011111001111111100011101000100011111111100110011110001111100000100110001000111111101000101010011011100110011010011,512'b01000000110111110111110100000111011100001101000101000011000100000001001111110001010001000100110101010001010001110111110111010100001101011111010111011111000000111111000001000101110000010011000011000000010011000011010101000111001101110100111100000011111100010100001111000101110001001111110000110011011100010101111100000001000001011101000001011100000101111101000011000111000101010001000111000000111101110001010111010000000000001100010011110000010101001111010011010011000100111101110000111111010100111111000101111111,512'b11010100001100010000010111010001010011010001110000010011010011111100110000111111110000001111010111111100110100000000000101000100011100000101110011000001010101011101011100110001011111000011110000001101000101111111000111110100011111010000111111110000000100000001000011110000000000000000110100111100000001010000010111001100011111110111001111000111000011000001011100111101010001000101111111110001000001110000000011000101000101000000011100011100110011000011000001110011010101110100000100000111011100010011001111000001,512'b01110001011101110100110001001111111100110000000001001100110111001100011111010011000000110000111101010101000011011100010100000011010011000011000001110001110000111111110111111101001101110111111100001100010100000000010100000000000101011100010100010011111100000001011111110001000101000011011101110001011111110111000000000011011101000100110101010011000101110101010000000011111111001100110000010000110000011100010001110011010001010101001101110100001100010101110011010101110001000100000000011100110001000001000000110001,512'b00010000110111110100011101010000110111001101000111110101110111111111001101111101010000000101010000111111010100000101111111001100000001011100010000000111010111000001011111111101000011111101011100000011010100110011110101110000110111010100011111010000110101010011010001110100010011011111011100010001000000110000000111000111110000000001111101001100010011000001110100110011110011000100011111010011110011010111110111110001110101000011010100001100011101011101000111110111010100010001000000001111001100011100110111011101,512'b11010101000111110101110000110000001101001101010101000100010011110001010000111111110001011101010001110001001111111111011111010011001111001101000111001111010100010000000001000101010100010001010000010100010101111100001100000000110100111101011111010011000011000101001111000100011111110101000001000011110011011100000100000011010111001100010000010111110100001100011100110011010011010100001100011101010000111111001100000101010100111100000000011111010001000101000111010101001100000011000101110111011100110100000001000100,512'b01010011010001011101001100001100111111110011000100010111010011001111010001001111001111110011010101011101000111010101001100010111110000011111110011011101010101001100000001011100010100110000110000110011000101000111000001010011001111010000000111010001110111110100111111010100001101001101111111001100000111111111001111000100000101110100000000011101000011000000010011110101110101011100001111001111111100000001010011010011010100001101001100011101010111010011011101111111010100110001110000010101110001000100111101010011,512'b11110001010111110111011100001101010001000101010011000101010011001100011100110100000001000000000101110000110011111101000011001111110111110001111100010011000111110111110001010001000111001101111101110000010011110100110101110011000011001101110111001111111100000100011101010001110011000011001101010101001111011111010111010111000001111100110101010101001100011101010000010001001111010001011101000001010011001100111111110111000100010011111101110001001100001100000111110000001100000100010000010011001101110100000001000001,512'b01110101000100010101110101000001010111010011111100010001000100001101010100000001110011110001010111001101010100010101000000010011110000010001010000110011110111110100011111010011000111110001010001010101001100010001110001011100001111000100010111010011000100111100000100001111110101110011010011010011001100010011010101001111111111000001000011010101010001001111110001110001010101010001110100010101111101111111110001111100010011000001000011110001010111010111110001011100010101010101000000001101000001010011011111000101,512'b00110100010100110000110000110011000000001101010101011111001100000100010111110100000100001111110000110011000000001101110000010111011111110000000011111100000101000001111101011100010000010111001100010011110011111100010000110101110100010100110011110000001101000000010000111101110101010000110001001111001100111100010000011101011100011101011101011101000000010000010001111111000111010001000100110000111101001100000101000001110011111100010001011100000100111111111101110111110001110111000111000100110001110101010000110101,512'b01000111011100010111000000000111000011001100010011001100011101001100110001111100000011000001000000000011010001000000010101000000010000000000111101000000000001001100111100110111110111110001010101001100011100111111010111001101011101010111010100000101010011001111110000110101000011010101111100001101000100010100011111110011011100000011110011010001011111110011000101110011000000000100011111000001010000011111000100111101011101001101000100000011111100000011010100000100001111011100000111111101010100010011110100110000,512'b11000000000111000001110100010011000001011111011101010101000000000011001101000000001100000011011100001100110001110011010101000001000001000011011101001100011111000001110100001100000011001111000000000000110001000011001111001111110011000001010111110101000101110100110000010111110101001101110001001100010001110000110101000100110100110001000011001100001101000000001101010100010001110100110111110111111100010000010111001111001100001111000001010111000011000001111100001100110100000011000111000001110111000111111100010101,512'b00011111111111001101110101011100010000010001111111110111111100110101011100000000110000110011000000000011011100011101110111110100110000010011000100010000010011010101111101010000010101001101000011000000010101001101011111010000111101010001000001110001011111110001110001110001010000111101111111111101010011011100111101001101110000000111000011010100010111110111010011000000110011000100010000001100011100111100110011010001000000111100010100001111111100010001110100000100010001000011011100001100010011000000010011001101,512'b01010001110100110101000100010101000101010011000101110111011111000100000100011100000001000001001100110001111100010111111101110011001100010100010111011100001100110111011111111111001100001101110101110001011111110101110011001111000000110001111100110000110001000100001100010011010101011111110000110101110111001111010111000000110111010001000001001100110001000101111100010001000000110101010100111111011100010101110011000001110011111101110001110000000000110011010000010111000000000000110100000001010111000001110001010011,512'b00010000110101000111110000000001010011000101011101001101011111110001000100010111010111010001110101110101000001000111000100010000111100010111110000000011010111110100010100011101111100010111000111000011110000001100110000010111000011011111010000001101110101010100010111000100110000011100010111011100110111001101011100110000000011110000000000110011001111111101011101110011110001010100110100110101001111110101010100011100110111000111000001110100000001001111000111110000110001000001110000010011010011010000000001000011,512'b00000000000000111111110001010111111111111111010001011101011100010001110111001101011100001100001101010001000000000011000001000111110000110101011100010001010000000100110001000001110100010101111100110100000111111101010101110111001111000001010011000111110111010111110100110001001100000111110101011100011111001100111111010000110100000000111101001111010000111101000111010101110000001111011100010111010000000011110100110011010000011101010011000000110011011101001111010001000001110011010000000001000001010000011101010011,512'b11001100111100010001000100111111110001111111000011011100010100110000010011001100000101000000110000011100010101010011001100011101001101000111111101011111010000010000000101001100010000001100000100011101010011111111010100000101011111110111110001111100000001110000110011010111001101000111010000010100111100111101010011111101010000000000010000000001001111000011000111011100110100010101110001010001001101000100110101000001010100001101001100000011000100001100000001000111000001010000110101000111000100110100110001010100,512'b00010001000001001101000101000000010011001101000001111101000111000001000111010011001111010011000101010011001100010100001111111101011111001100111111010100000101010001000000010100000001000000011101010101010111011101110001011111110000011100010011000101111101000001110011110100110100110101011101011100110000111100011111001111010000010100110000000100000100001100111100010111001100000101001100010000110101000101010001110000001111110011000000010011010000001111010111000000001101010011110100110111111101110000000100011100,512'b01011100110101010001000100111111001111011101010100001101000100110100110111000001111111011101010000000111111101010100000000000101011100110111110011110100000111010111010111001111000111010111110101001101110101000101011100000100111100011100010111110100010101010100110100010000111111000100111100110001111111010011110011111111111101111111110111011100110000011100001100110111000111000101110100001111000111000111011100001100010100000100001101110100010100000111110100000001001111010011001111110000110011001111001111001101,512'b01110100010101010111001101011111110001000011110111110000010011110111111100111101000000010000110101001100111101110001001111010011110100001111000000010000000100110101001100000001000100001101110001110111011101111101000001010111011111110001000011000000010101011111010011011100010101001111001111110100010111111111000000000111000000010000000000010000000100000011010011110000001100000001001111111101001111001101110001011100001100000001011111000000110100011111010000110100000011010100010100001101110011010101010001000011,512'b00000000000011111111110011010100110101001111111111010100001101000100110000010000110001110101110001111111110111001111000111000000110000001100010011000001000100000101010101001100001100011100010111000101010000010001010000011111011101111100000000111101000000010100111101000011001100011100000011010100010111110101010000011111110011011111000101000100001100011100010000000111010111010001001111010100110001000000000000110100000011000100010000000000111100110011000101110111001100110101010000110100110000000000000101001101,512'b00010000000000001100000001010000110000000001010011000001000000011100000001010000011111000100000000000000011100010001001100111100010001110111110101110011001111111100010111110101000101110011000000000111110100011101110111110000111101110011001100110111001100001101010001001111000100000011111100111111110111110000010011010100000001000111010100010000000111001101000001010101111101110001010111010111010000011101110101010111010100000001110000111111000101010101010111110001110000010111001100000011110011110000010101011111,512'b00010001000001000111110101000100000100110011011101001111011101010111001101010001110101001100010101000101001101000100110011000011001101110001011101000111010100000111000101110100001101000000110000110100000011010011000111110000000001000001110011010001000011010011111111000000010101001100000000011100000100111101110000110011000100110111000100111111001101110001000001010000000011000000001100111100111101011101010001000111011100001111110001011111000000001100001101001100110100010011110111011100010001000100000100010001,512'b00010011001100010100011101000111000001011111001100111100111101110101000100010011010011010111010000000000110111010001010001001100001101000011110100111111001101110101010001001111000000001101010011000011110011000101000011001101110000111100111100010000111101000100010011110111111101110000111101111111111100010100000111010000010111110100001101011101010011111111010001001101001100011101000101010111011111011101010111110100000111110001000100110011110011000100000001110001010100000000110101001100001101010011110111001111,512'b01000001010100000000000111000011010001000101001100111101000000110101011100110100110100001111000000000101001100010111111100110001010100001111000001010000111100000101110001111111110100000111110101001101010000110001000011111101110101000101110000001111001100001111000011000111000001110000110101000101001101011100001111001101010001001101111100011101110101111101000001000101011100111111010100001101110000111100011101110000010001110111011100000001110011000101000100010100011100010011000001110100111100011111010000010100,512'b01110000010101011100110101010111111101111100010011000001011101110000010011110111010011000101110000110000000000001111110011010011000000010001110011000001000111000100000100010000000100000101000100011101000011001111000001010011010000001100010011110100010011110001000111000001000011010111001100000000000011110111000001000001110111010111110111000100010001011100010111111101011100010100000111000111000111110100111111011101000101011100000000010111011100011101000111001101110000001111000000000100110100010100010011000111,512'b11000011000111110000010101111100011100001101000011000100011101110100010101011101001101000011010111010000001100000000011111110001000101011101011100000000110011000001010111010011110101011100010000001111011100001101110100110011110000110001000100010100111101000101011101110100110101010001110011110011110101011101010111011111001101111111011111110100010101010000000000110101111101110011011101010000110001110101000011000000001101011100010111011111111111111101000001000100001111010101000000011101010100110000000111000000,512'b11000101010101001100010011001111111101000101010001110000110111000011000111010001010001010101111100001100000011110011110000011101111101001111110111000000110000000000110000010000010101110000000100010111001100010101001100001111000011000100010001011101111111001101000100111101010001011101001101000101010000011101011111001101011101010101001101010101000101010101111100010111000000110111110000000100000100000001000000110000010100000101010001001101111101000100000111111101110011110111000000110000000111011100110001111101,512'b11010011001101111101010100011111010000001100010111111111110101001111011100001100000100110001001111000011010100111101110000010000111101000000000011111100110101110111000011110101011111110111001111000011000001011100000100111111110111110111001111011100000000111100011111000011010100010001011111010001010111000100110101001111010100111101111100010011010101111101001100110101010100110001001100010111010011000100110001111111110100010000111100011100010000111101011111110100111100110000110000000100110111110101001100000011,512'b00000001110101111101111111010001001101110100010011000100110000110000001111010101010011110111110100110000110101001100111100000111010000110101000001000001001100111100110011110101001100000001111101110100110100000100000000110001000111001100001101111101011101000100000000000001010111111101001100001101000011010100111100010001000100110011000100000000000100110011001100011100011101011100001100001111000000000111000111110111010100000101001111010000110001001100000011110100001111110001010000000011000100010001010001111101,512'b01011111000100000011010000000000011101110001110000110000010111000000011101010100010001010000000100001101110000011101001111110101110101000100010111111101010111110111110000001100001100000000000001110000000100110101111111010101000100110000001100000001010000010111000000110111110011110001001111010011010001110000110000010000110011000000000011110000000101001100110111000101010100110111110001110001001101010101011100010000010011011111000001111100010011110111011101000000001111001100000011110100010011011111010011011101,512'b00000101110100001111001100000100001111011111011100110011110100010100000011000100000101000011011101011101000011000100000011000100001101001101010011010000110100000011110101010101011101010100001100000100111100110011110011111100110001000100000011010011001101010011110100010001010011000000110011011101111101010011000011110011001100000001000011010101110001010001010111010000000101011100001111000000000011010000010100011101000111110001110100010001000011001111111100110100000001000101011111000000110000000011010001110101,512'b11110100011100010000000001111100011111110100000000001101010011111111010101000000000101010001000001110100011101000100011100001100110000111111111101111101010001000100111101000001111111000111010111001111010001010100110000010101001111011111010100011100011100010000010011110001001101110000010100000011011100000000001111010001110111011111010000011100011100001101110100000101000001110000001100110111000000000000000100001100001100010000111100011111010111011100110101010000110001011101010011000111110000011100011100000101,512'b01000011111100000111010100001100011101000000010100111100000111010000010001000000000000011100001100110001000111111111011111001100010001010111010011010001000111110101110100000000011101010111011111110000000001000100110101010011110000110111010111000101000111010001001101001101110011001111110000001111001111110011000011001100110100111101010101111111010111111111000101000011010100110100110101010100110100001101000101110100000001110000010100001100110011010000011111111100110100010000000101010011010000001100011100110000,512'b11110011010100010111001100010001000001001100010100010100000001010000110111111100000100000111000011001100110111010001110001110001010000110100010001000100111101110101110111000001000000001100111111001100011101110111001100110011110011111101000111010011000001000100000101010111000001000011011111001111000000110000011111001111000101001101000000011101110000010101010111010000110100001101110101010000110011000101001100010011000001011100001111000111011101010001110101110001000000000100110100000001010000000000110101110001,512'b01010111011100111101010000111100000001010101011100001111111100001111010111010011011111000100111111000100000001000100111111000101011100111111110001001100001100010000011111111101010001001111110100000111010011000100110100010100110000000011000011010001110100000001110000001111111101000000111101000011110000000000011100000100010111110100010000000111000111010011010100000111001111010000110001110001000111010111010000010100110000000000011100110001000011000100110001000000110001011111001100000000000101000000000001010000,512'b01000011000001001111010000010111110001010001010001000111111100010000110111000011010000110111000011110000001101001100010100000111000000000011110011111111110000110001001100010000000100110001110100010100010101001111110011010101001100000100000000000100010001000000110101001101010000010000110001110101010000011101000101110100010100110101000001010101010111001101011111000100111111110011011111111100110011000111001111110101001101011111110011001101011101010000000100000111010001110100111100110100010100010000010011110001,512'b00000011011101110100001101010111110111111101010101110001110011111100010101001100011111001100110001111101010101011101111100000111001101011101011101111111111100010100000000000011010001000111111101001100110011110101001111110100111101001111010101010100111111000101011111010111010000010000000000110001001101110100110011011111010101010100010001010000001101110011011101110000000100110111000000001101011100000000111100011111111101110101011100110101010101010001000001111101000001000111010000010011010111110011011100011101,512'b01110101001111000100010000001101010001001111110000000111001101010000010100010101011100010011001111010000110011010011000100111101010101000000010000110111000000010011001101000011010000110000001100011101000111011111000011111101001101010001111101111100111101010101001101000000111100000011000001111101010000000100110000010011000011000101001101000011000111110101010111110111010100010011010111010011110001000101000000000100110011110011011100110101001100011100010001010011110100001101000101111100011100010011010000010000,512'b11000001000000110111010000111111010001110100000000010000000111011101010001000100000100010100000001001101011100001100110000110001000000000111110001110100000101001100001101110101111100010011001101001111110011110011110111110100010011110101110101111111000100110001110000010111010000110001110001110100000011000101000011110000011100010100000101010100000011010111000001010111000100010101110101000000000000110011010000010001000001000111010011011111001101000111010011010100001100110101010100110100000111000011000001110011,512'b00011111011101010111011111110101011100000011000100001111001100010100110001000000000011110111111100110011000011001100000101010100111101010111010000001100000101010000000111001101111100010100110000010011001111001100110001000100001111010001110011110100010011010111111100000100001111111101001100010000001100001111001100011100111101111100111100111111010001011101000011010111110011001101011100110111010100010100110011010101001111000100001101110111000111011111010000010000111100000000010000001111110111111111000101110011,512'b11010101000011000111110011000011010001001100111100110001000101000000000011000101001100110011000100110001011100010011001111110011000111110001001101000100110100000011001111000011010111110000001100010001000000011101110001110000001111111101000011110011001111110000010001001100001101001101110000010000010000001100010100111101011100010011011111011111001111010000000101110001111111110111111100000011010000010111010111110001111100010011001101110000000111000011010000000000010100000001011111111111110100011101110101110011,512'b01010000010011010100010000000001010111000100011101111100110011001100110101001100110101010011111111010000011111011101000000111111010111110001010000001101110101010001000111011101010100000001000000000111011101011101010101001100111111001100010011001111110001110011110101010100001101111101000101001111000111011111111100110000000011001100000100000000000100110000110001001111010101111111111101110001011111010011110000000100010101010011110101011100110100110000110011111100110000110101010011110001110111111100111101001100,512'b00110100110001110100011100001100010011010100110101010100001111110111110001010100010011000111110011000001110001001100110011010100001101010100110000001101010101000100000011111111000000111100110001011111110000001101011100000011110001110000010001000000110011111111010101000000000111000111010000000001000100010100001100110000110111000101000100110000010000001100000011110011001100011111000000110001001101000101110111000100000011110001000001011100110001001101111100111101110101110001010000111101110011110000000000000001,512'b00110011010011010000110111010001010100010011000101111111000001001101110100011101110011001101011111000100001101001101000001011111110001001101010000110111111101010001111100111100010000010101110000011111000100000111001101111100000111010000011111000000111111001100000000110000111111110100010011001100010000000111110000111100110000001100000111110101000001111111000011111100001100010011010001000000110100110100000000000001011100000011110000010101000011110011110101010111111100001101010111011101110000011101001101000111,512'b11111100111101010000011100001111010000000001001100010101110000000000011101000001111101110011010100000001000101110000010011011100000000111111110001110011001100000000000111111100110000110100001101010100000111011111110011011111000001110001011100110101111111001100000111110001000100110111111100001111010100010101001111010011000001000011000000110011001100110000111101000000011111011100000001011100000111110111111100000100110000011101000101010011011100110011110011110000000000001101110111011101110000111101110111010001,512'b00010011110111110001110111000001000000110101011111110001010100110100011100010000111100110101011101010000110011010001001111000011001101010000010111000100010111111111000000000011110101000011001101110001010101001111000000000101000000001111000100110100000000010000001111010100110011000111000100010011001101010000000001000000001111000100000011010101001101011100001111010001010100001100000100110101011111001100010111110101000111110000000011011111110011010000111100110001000001011100010001000011000100010100001100000001,512'b00000001000011001111000100001111010011010000111111110000010000110001010111001100010011000001111100110111010101010001001101001100010000000101010000010011000000010000110000000101111100000101000000001101011100000001001100111111001100010101001111000000110111000100111101110100001101001111010001111111000000001111000001010100111101011100010000011100001101110011110101110011010101110001000000000011011100000000000101110100010101011101001101111111111100110011000000000011000101110100010000000000111100010101010111000101,512'b00010101001101001101010100111101011101110000000101000111000111010011110000010111010000110001001111010101110000010111011111001100000000000000010101010111110101011111010101000000110000010100111101001101000000000011001100001100000001000111110111000001111111110101010000110011000000001100010000011100010001110011000011000101111111110011110001001101010111010001010111111100000000000011010111111101001101011100000100010011010000000001110000011101000000110111001100010100110000001100011101000000110011110101000000110000,512'b00110011110101010100010000001111010011000000001101001111001111010000110000010001000111110011111111000100000100110011000001110011011111011111010011011100000001010111010001001100110011111100110011000111111101000100111101011101110011001100010101000001011100001101010011010100010100010101110001111100011111000101011100000011110001111111111111001101010100000001001101000000110111000000001111010101001101010111110000000001000100011100111111000011110111111111010001010101110000010100000000001100000101011101001111000001,512'b11000000011111110011011111010001111111010001110000110000011101011111000000000011000100111111011101000011000101110000111111011101011100110101001100010100110000000001001111010111010100111100000111010011010101110111001111110100110011010111110100111100011101000000000111001101010011010100000011001111000111111111110001001111000000110101110100000011110100000100110101010000110011010111110000010000000000110011001100110011111100110100010001111100000100110011001111110001001100000111110111010000000111001111111100010000,512'b11000001000111000100000001010011000100010001111100110001010100110001110101010001111111000000000011010001000100110101010111110001000011000011110101010100010001111101000011110101010111110000110100011101110111000100110001110000001111111101110000000001111100110101001101011101010011010111001101110100000101010000000000001101011100000100000000011111010000110101000001000001000011110001000101010000000111110000000000010100011111110011110000000001000011000011001111010100000101000011000100000100011111111101000111000001,512'b00011100110001110111000000000000110001111101000101000001000111001100010011000100010000000111010100001101001100000011000000011101000011111100011111011101010011110100010011000101110000000111001100000111110000001111010001011100110001000011001100000000010111010011011101000001010001000111000001000111011111010100011111110100010111000101110001110001010000000100000000011101111101000101011100110000000001111111000100010001000101110011010000001111001111000000110000000011010111000100010001000000010100110011011101010101,512'b11011111111100111100001100000111000101011111000011001111010011110001010000110111011111011101011100011111001101001111000000111100010011010011010111110011000100110011000011110100010001000100001111001111000000110001001100000100001101000100001100000111111101001101010000000011000111110100010101010011001111010101011111110000000100110001000001111111000101110101001111000000110101000000000101011111111111000001010111010100000000000000000111010001000100010100110100010001110101011101001111010011110000010100010001000111,512'b00110011001100010011010100000011110101010011110101001111010101010001011101010000110000110011111111110100110000010001000001011100010000110001110000110000001101011100010011000000000000010011010100010000011111110011000011010011010111011101010000001111010111000100000101111101110000000000110000000100010101010100010000110111010001011111111111000001000011000011010100000011110111000111011100010100000000011101000111010100110001000011110000010111001101011100010101011100110111000100010000010011111111110000000101111100,512'b01111100011101010011010001111111111100110000011101010101010101110011110100010111110101011101000101010100011111001101010100010011110000000100001100011111010000110001010111000100000101111100010100111111000101011101010111000101111100010001010111011111000100111100010001010001010011010000111100001101001100110100000100000001110101001101110111010000011101000001010001110001110000000101111101010001001111000111000101000111110111010011110101110100000001110100000000000011010011001101011101011111110111000111000011000100,512'b11110100010101010111011111010000111100110111010001010001001100000000010100011101010000011101110111010111011101111100011101111100000100110011110001000000000101001101000011110001011100010001000001010111010011010100010111010000011100000000110100110011110000000100111100110011000001000011110001010000001100110101001100001100110100010000110101010000010100110000010001010000111101110001010001000100000011111100010000010001110000110000000011000000110101111111110000011100000100011111001111010000011101110011110011000001,512'b00000011010101010111010000001100011101110000011100000111000011010011000001000100010000010000001111010100011100110101110101010011001101111100001100011101000111110101110111001101000011000011010000111101001111110000010101001100111101000011000011000011011100111100110000001111000011001101001111010111000011011100001101000101111101000001000001111100000000011101110100110111011100011111000100010011010001110111000111000101001100110000010001000001000100000011010011110101110011000011011100110101110100000000000100010100,512'b01000100000011111101010100001111110101110100001111110011000011110001001100110101000101111111010100000001011111000000010100010101010000010001000011010011110111001100110011111100000000010000011101001101000001011100000011011101001111000001011111001100110100010100000000010000001100011100110000000101010001000000001111000101010111010100010011110011011100110101010001110001011101010111110000110111010000010001000111001100010100111111011100010001000100111100000100011100010101111100110000010011001100010000011100000111,512'b11010011110000010100111111000111111111111101110101011111000011010001000001001111000101000011011111110101010100010011001100011100010100001100110001001101000100011100000001111101111100000001111111000000000011001111110000001111000011000101010001111100111111000101010001001111000000000100011101001111001101000100000101110100000111000100011101010000010001000001110011001100110000111100110001010111111111000100000001010111111101001101010000011100110111010111000101110011110011011111000011011101110011011111000011000000,512'b11000111000001111111110100110011001111000000111100001100111111111101110101110101111101011100001101010011000000010000000111110000111101011101110101110101110000000000000011010100111100011100000101110011010011000011010001010100010000010100010111001111111101110101001100110111010001010100011100110011110111000100000101110100000011011111111100000100001100110100010100010100110001000001010001000000111111110011010100010101000011001100010000000011000011001100000000110101010011000111000000011111010101110011110101110001,512'b00001111001101110001001100111111110101110100010001001100111101110111110000011101000000110000010100010001111100000111110111110000000001110100000000010100011101010100011111000011010001010001001111000000000100000000011111011111011100000011011101010101000000000100111100010000000100110111001111000001001100000101110001110001110000110001111100001100010000110000110101011101110111000000011100000101011111011100010100000000000000011111000011011111010011010101000100010000010000000111010011010111110000110000110000010000,512'b01010000010101000100010101010011110011110100000000110001010001110001011100000100010100011101010101000011000101110000000000001101000011001111110111001101110011110000110000111111110011010000010101010000111101110000001111000000110001000111111100010000110101110001000000110001010000010000000111110111011100110101010100110000111111000100010001011100010000011100000100001101010111110101011100001101011111110001000001010111001100000001001100000011001100110000110101111111110011110000111100110001010000010111011111011101,512'b01000101110111000100011111001101010011000111010011010000000101000000001111010111110001110001000000110000000000110001010001001111110011011111010111110000011101000000111100000001000001000001010011010001010100010100000011110011000100001101000100010111010101000011110101011100010000011100000100000101110100010001010000110011010100001101001111110100000011111111010001010111010101000001111111010111110011010111010100001111010001111100110000010000000101010101111111011101010001010100010011110100110111110011000001000100,512'b00011101010111110100001101011101010011000011000101010101111100001111010000110100110011000000110011110111010000010000010111001111010000110101110000110111110101000100000011000001110011000100001101010000110101000100110101111101000001111101110001110101011100010100000111001100110011110000110101000001000100011101010101010101111101000111110111111100011100110100110011110011010011110001001101000001001101000001000011110011010101000000010101110011111100010111001111110100110000001100111111110111001111001111010100011100,512'b01110001000101000011000011010000000011010111010100000101110000011101010000001100000000000000000001010111000100110001010011000001000011001100111111110101000000011101000100010001000011011100000000010000010100001111110111010111110001010011000000011101000100000100000001011111000000001111001100110111000001011111010111110001000111011100000011011100010111111101111100001111110000000000111111001111011111110000000011110100001111000000010100110000010001110111001111111111010101010000001100001100111111111100010100010011,512'b00001111001111010011000101110011110001000011000100010111110111000101000111110001011101110001010111000001011101011100010100000001110101000011011100010000110001111100001100000111000000111111010111110011010000000000110101010001001100000000110100001100000101000011011100000000110100111111110000000001011101001100010011111100000100111100111101110000110001010001000000011111110000010100000001001111110011111111000101001100000011000000000100011111010011010100011111001111111100010000110100010100111100011100001111010100,512'b11010100001100010011000111001111110111001111110000110000000011010111011101010100110100000011011101110101111101000111001100010111011100110011110001001100111100110101000011001100110001010011110000110000111111001101010011001111000000001111000111000100010011000001011111001111000100000111111111000011110001000001000000000100001100001100111101000111110111010001010100010011110100010011011111011101000001110000010100000101110001001100010001000101000111110000010100110011000111011101010101111111000101010100000111011100,512'b11000101010111001111000101000011011100010101001100110000000011010000001111001111001111011111110011000111000100111101000001110011000101000001000100000101010000010011011111000101111101110111110000000000110111001100000001110111010101000011000001111101001100110011011100110001010001000011111111000000010111011101110001010000000100010100000111010000010000110100000101011101011100110111010000011111000111000011111100010000110001000100001100110001000100110000001100000000110011110101111101110100011100010001010101111101,512'b00001101000100011111110101111111110101010000110011110111010111110001110011010001000011010100010011111111011101111111110000110111110100010000001111000000111100000111010001001100001100011100110101010111011101001100010100000101110101010001110101110000011100111111000011001100000011011111111101110101110101000001111111110000001111110101001111000011110111000111010100001100110111110111111101011101010000011101110101010101111100110011110100110001010011011101010011110001000111000000111101010001111101110000011101000001,512'b01000101000111010101110000011101110001110101011111010000111111011100000101010101110000000001000100011101000100010111000100001100010000001100110000010101000001110100010000110000001100110000000011110000000111110001110000010011111100010111001111010100011111011111010001000011010100000101000101010101010111111111000101000001010101010011000011011100010111000111000001110000000000011111001111000011011101110001011100001100010011110011010100011101000000000111001111000111011111010001010100110100010001000101000100010111,512'b00010100000000000111000100001100010101110001111100010000110101010100011101000011010000000001000101110000010100010000111101110001010000111111000000111101000001000011010100001100011111110011010101000101000011110101001100010011011100000111000111000001111100110011010011010001000001011101010000000001010000011111000100010111110101000000000100000011111100010001110100111111110100000000010011110101011111011111000111011111010011110101011100110101111111110001000111001100000001010100110101110101000000000000010100110000,512'b00111100000111010100010011010011001100010011010000000000011100000101110011010111111101010011110000011111000111110111011111011111111111001100011111010001000000111111000111110101011100001100010100111111111111110101110001001101011100010001011101000111010001010000000100010111010001011100001101010000000001110000110111000101000001110000010011000001001111000101000000111100000100010100011111001111010101111100110000010111111101111100000000000111010001000001011111111101011111110100011111110100110111010101000111110001,512'b11011101110101010011011101001111000000110101000001010000111111001100001100010001000101010001010101011100000000011101110111010100010000110000011111000101110001010011110100111111000100001111000001000111001100001100010000001101000111011100110111010000011111001101110011110100001111001101110011000000110001000100110111010011001101001111001111110000110111001111110001111101111100001100110001000000010100000000000011110100001111010000001100000101110001110000110000001111011100000101000111010100010000111100001100011101,512'b00001100000100110011000000000001011101011111011111110000000000010011001111110000110001000000000100111100110101010000000011110111010101010101000100110101000101110100010011110100010001000100110100110001110011011101010000010000011100110000110011010111010101011101000011111100110001000011010011011100010001111101110001001101110000111101000011110001001111011100000000000001011100000100110101110000110000010000010000000011110111000101000111001101010000000000111111000001111101110111010100110100010000011101000111110100,512'b00000111110100110111111100000011001101001101001101110111110001110100000000110100001101010101010000001111000001010101000001000100000100001101000100011111110111000001001100111111110001110011000000001100001101111100000111001100010100110111000111011101110000010101111101011101000011000000000000000100011111010000000001001100000111000001010101111101001111010001010100000000010101111111010111000000011101001100110011001111000111000011011100010011000100001100111111110100010100000001111100010001010000110100000001010101,512'b00010000010000001100111100000011000011001100001100001111000101011100011111010101000000011100110011110001111101000001110001110101010101010111111100010011000011110000000011000001011111001100000001111101000111000001010111110111000011000101110111011100001100011101111101001100011100110011000101111111111100110111010111011100111101010000001101010101110111110011000011010101000111001101000011000101000111000100111111110011110000110000110000000000010000001111010001111100001101000101000101011111000000110011000011000100,512'b00001111010101110011000011000100010000000100011101000101010000111111000101110100010001010111011100000000001100010011010000000100001111111101000011010011000101110001001100001100011100011111010100110000110001110100110011000001010100010100000001000011001100110101110011010111110101010001000100001100000011010001110001111100000100001101011101111101011111110101110000011100000001011101110011010100110101000100010101011111011101110000011100010101110111110001000101001100000100110000110001111101000001000111000100110011,512'b11000011010100010101000100111101001101000000011101000000000011000101010000000111111100111100010101001101000100111101110101110100110100001101010001000100110001110111111100110100001111110100010111111100110001110001111100000111010101010001010000010101011111010011010000000111010100110001110100011100010000000001110100010001001111011100010011001100010000111100111111000111001101010100000001110011110001111100011100111111010000111101001111111111110111010011000011110001010011001100111111011111000001001101011101011101,512'b11110100010111000000001100000000000001001111111101000111001111000100010111110001110001110101000101010100010000110100001101000101010000000111011111110001000101000100010000001100010111000011010011000000000100111111001111011100000111000011000001000001001111010100000111010101111101011100000101111100111100010000001101000100000101000000110111001100000000010011110000011111010011011111001100001100011100110011111100010100111101010001010100111101110000110001000100000000000100010000000100111100110000011101001101000011,512'b00001101110000111111000101110001011111010000001111010101000000000101000000010111001100000101111111000111110001111100011111000101000000110011111101111111000000011111011100110001010001011101011100110011000100110111010100010101001100110000000100011101110100001101000001111100010011110001000000011101010111010011010001010100110011000000001111111100010001111101011100010011110011111100110111011101011100000111111100111100110100010111011111010111000001110000001111110101010000000011010101000000000000001100010011001100,512'b00111101110111110011010000011101011101110101010100001100110100001111011101111111001111110001000101000011000100011111110111000000010000000000010011000100000011010101010001010101110011001100000000011100010011110111000111111100010111000100000111000101110111011100010101110011110100000000000100010100111111001101010000000000110101001111010101111111000100001101011111010111001111111100110101001101010000000100000001000011010011110101011111010111000000000011110001010100111111010011000001000100010000110111000000000011,512'b00010100001111000111000001000100000011111100011101111101111100010001010011000101010100001101110000011111000101010011111100110001110001000011000000111111010000000101000000001100000001000101010001000101000100000000000011010100000011000001001100011111000111111111110000000101110001010011011111111111010101111111110001001111000100001100010100010000110011000100110001000000110000000111010011000000000001110000001100111111000111010001000111110101000001010101001111000011000011010100001111110011011100111100110011111111,512'b11010100010001010000000100000001111111110100010000001101011100011100110001111111110011001100010111111100110001011101000000110001001111000101011100110001011100010001111100110011110111011111000011111111111101011111010100000011000101110111010011001111001100001100000000110000001100010100000111000011011111000001110111111100000100011101000000001111000111010000110000110001000101011111010101010111111100110101000111000011000100000000010111110101110100011100001100010000111101010100010100001111010111010111110111010100,512'b11010111000111011111111100001100000100111101111101000000010000001101001111011111110100000011000001000101001111011111000000001111010011010000110000000100010101000011010001001111110001001100000001110000001111110100000000110101110001010011001111110100000000010111011111000111111100010000000100010111011111001111000101010101000000111111011111110000110100001100010011110001110001010011000011000100000100000011000100111111010111110000010111010111111100001101010111111100000111010111110101111111111100000011011111001101,512'b11000100000011010000000001001100110100110011011100111111000101111101000000111100000000000100010100110011110001000111110001010000110111110101001101000111000101110001000100010111001101011111111101110001000000010011011111001101110000001111000000010001010000010000000011011101000101010100110001010101010000010111011100110000010000010111001111111111011100000000110011000001010001010001000000001101001111000000001100000001010101011100000111001111000101011111111111010001111111000111111111000100110000001111110101000000,512'b00010011110011000111001101011101000100110000001100110001001101011111000101000001010011110111010100010001011100000111000001110001110000110001000000010001000000000101011111011111000101010100011100001111111111010111000111110000111111110100000111000001111101011111010100110001000111110111111100011101001111110111010100000011011111110111000101000100110111010100011101001111010000000000010100001100011101010111111101001101010100000011110011110000010111000100110101000011110100001101000011000111110111111111000000000000,512'b01011101000001010000110000001100010100110100010001111111001101110001001111010001000000011111010111000001111100000000110100000000110100110111000001110101111111110001110111110000001111011101010100110111000101001100000101010011000011010011110100111101111101001111001101001111110011110101001100010000001111010001010100001111001100000000001111000011000100001111000100111100011111000011110101001111011100011100000111000111000011001111011100000000110101010000000111011100010111010011001100000001000011011111011100111111,512'b11000000000100010011110100110000000011000111110000000011110000111100011100000101010100000101111101000100001111110000000011010001001111110011110000010000111111001100001111011101000000000000001101000011010111000001001111000011110000111111001101110101000000000100001101011100001111000111011100110100110011000101011101110001010100110001001100000011111101011111111101000101001100010101000111000100010011011101011101001101010101111100000101011100000000001111110111001101010000110101001101010101110111010101010101110000,512'b01000001001101000001010011001101000000000111011111000011000011000101110101010100001111110101000101010101010100000000010000110100000111110100111101000001001101110000001101011100000111000101111100010000110011001100110111111111111111000011000111110000011101010101010111001101111111001100110100001100000101000000000001000100000001011100110111000011111100110100010101000001000001000001110100010100000000011101010011010100000000111101000111000111110100010001000001000000000011001100000001010100111101011100011100011111,512'b11110111010011110000000100001100011100011111011100000100001101011101010101010011000000001111011111111100011100001100011111010100110100000111110101110011000000000111001100000100001100000111110100000001000000011100001111111111110101111111010111111100000111000000000101001111000100011101110100000011010100001100011101011101110011001100111111000111110000001101110001011111001101010101001111010111000101000000110000011100000011110011110101011101111101111100000000000001111100011111010000010001010100000000010011110111,512'b00000011110011111101011101000111110001011101001111110100000001001100000100011101111111110000110001000101001111000011011111110001010100010011001100000000010011000100010100111111010101000111011100110001110001110101001101000100000011000000010000000001110001010101000101010111010000000001010000010000111111000001001111010101111111110001010100111111000101000011010001010011011111001101010011000111010100000101011100010011000111111111000101010101110100111111001101111101000100110100000001000001011101010001111101010001,512'b11110100010100000000000111000100001100001101010101010000000000000011000111110011110111001111010001110011010011001100110111000101111101000101111100111111000000010100110001001101000000000111001101110011010111000000010001001100000100000000110101001101011111010101000000011101000011000011010001000011000101001100011100111100000001110101001101110100000101000011110001011100000001000100010001111111000100110011000111110000110111000000000111111100000011000111000100001100110111110001000000000001110111010001010100000111,512'b11000111001100010011110000010101000001110101010100000000011100110000000100111100010000000000010100001111111111011111010111010101000101000101000000000000010101011101001111011101010011010111110001011101000011000000011101111111001101110101001101111100001101010011000011000000010000000100111111110011000001000000000101010011111101110100010101111111000111110000001111010001010100110000000101010001111101011101110111010000000001011111010011010100010111011100011101000111111100110100111100111100110000000100111100000100,512'b01000100000000000001001111110111001101011111011101000001011101111101011100011100000111000100001101011100110100010000000011010100111101001101110000000111110101110001000101001111010000110111110001001100110100111100110100110000110100000011110100000011001100000011000100010100110000000011110011110111000001001101110111010001000101110000010111000011001101010011000011110001010111010100000011010000000100010100000101110011000000111111000000010001011100000000010001110000001100000101111100000001111111001100000000000100,512'b11010000000111010000001111110000010101010000000111000100010100010001000000110011000101111100010001001101000101000111010011110000001111000011001100011100110111011111111101110011010111000001110101011101010101010101011100010000011100011100010000010111010001000101111111010101000001010111011111010100010100000001000100000100010011011101001101111111000111111101000000110001110011110001000100011100011100000001110001111111110001001111001111010011001101010100111101010001000100000001110000000011110000001100000101001111,512'b00000011110101110000000000000100001100111111000000110001010111011111111111011111001100010111010001011101010000010001001101110100110001011101010011001100000111000101110011011100111100110011000000111111001100001100110000011101010011110000010000010001011101110100001111000001011100011111010000110111000111110111110000000000111101000011010000001111010000001100110100001100110101000100001111000100000111010100001111000001010011010111000111001101000101110011001111110100010000000000110111001100110100011111011111110100,512'b11010100011100000000111101111100001111010111001100111101110100000111010000110001001111000100001100110111000111111111010000110101110000111111001101110001001100000101010001000101010000111101010100110100111100010100001100111100110011111101000111110111000001010011001111111101010111001111000000111101110101110101010101011111000000010000000111000001000000111100111100111101011101000100111100000100000000000111110100011111010111111100010001111101000111000000111111010111010001001111010011111100000111111111110111110000,512'b00000100010001010001111100011100010100000001010111111101110001011100110111110111110001001100001100000100110100000100001111011101010000110000010000000011110011001100000001110111110101011111110101010001001100010111000000110011001101011100000111001111010100111101111101001111000001110000110011000000111111000001011100000001111100001111110100111101011111001100000100000101011111111111011101010101111111000001111100011111110101110100000111011111110111000000011111110001001100110000010100111111001101001100010111000000,512'b00010100111100110011000001000011110000000000110111011100110101110000110101011111011100001111111111001101010111111101001101010011110100000001110000011101010100111111010000000000010100011100110100000011010100010100010101111111000101110001000011000011010100000111110000001101000101110000110100010100001100110000010111000001110101111111011111010000110111110000011100011111000011111111000100000000000111010100111101001111111101000001010000000011010000110001010000010011110000110001001100000011000000110000110011111100,512'b00110101010111110101010111110101000111010000010011010000010111010101110111000100010011001100010000000100001100110000110101000001110001011101110011110001000000000101110100001100011111000001000000000000011100011111000011000000000111111101110100111101000000000011010011000101110001000000111101001111000100000000011100111111111101011100000100000101000001010001110001110000110000000011010111001111111101110101110100111101010101001101000101000000001101111101010111000101110011000000000101010101111100010101001100010100,512'b01000000010100111101000001111100000011000011010000001101000001110001000111111100000101000000111101111111110101000001110000011111001111000100010101000100000000000111000011000011001111110101000001010100001100011100011100010100110000011101111100110101000011111101010000010100011101011100000100001111110100000000010011011101000000010001111101010001000011011111010111001100111111000000010111000100001101110101000000010001110011001100110011110101110011000011001100000001000001010111000100001101011111010100001101000101,512'b01010100000001110000000001000001011100010111111100001101010101000001000100011111111111110011011111000100000011110100110101010111010001110000010101010111110001110000110001001111000011000011110000001100111111001111010001111100001111001111010011111101000011010100010100000101110111000111011100010001000001011101111101000100110011000100010101110000000111011111110001010100110100011100010011110000010111111101010100001100001111000101110001001100001101001101010100011101110000111111010011000101000000000000010011110100,512'b11010111010000011100010100000000110000011100110000111100010000000100001100010000110101011100110000000001010001001101011100000001110000001100001101000101011111000101110101111111010011011111010001111100000001111100110101000011000111000001000001011100110011011100111100001111000001010101000011010111010100010101000111110011011111000001001111010000010000000001010000110011000001000011110100001101000011000000000101110000110101010001110000001100010111000100000111000101110101111100010100000111110000010011011100000101,512'b00110000110000000000110001000101011111110011110100010011010000001111000001011111010101010100010100111111110100001100010000110100000000001101110100011111110011110100000011000000010101010100110100011101011100001100010000110100110000001101000111000101001111011111110000010001000000000111010001110001110000010100111111110011001100010001110001010001110100000111110001000000001101010111000100010001011101110100110011110011111101001101000000010000000101000011001111001111000101111100001100111100110100001111011100010111,512'b01111101000001010000111111110100000101110001110000110000111111001101111101001101000000000111110101110101010011001100110101110001000101000000001100010101001101001100110000110100000011110111010000001111000101000100001100010111010011010101010001000100000000111101111111000001010111011101111111110100010001000001001100001111110000110101000100110100010000010101001111000000110011001101111101000111011101111100010111110111001100000011001100110001111111000011000101001101000011010000010000001100000001110000000111000001,512'b01011111000100000100111101000000110101010000000001000111010101001100000001000100110000110111001101010100111101010001010000110011000011110000001111111100001100010001010000010000111100110000000100010001011101010111110101010000000100110001000011010101001100111111000001000001000111010001000011010011010000011100110000000000000011000011000100110001001100000111000000000001000100001100000001010000110111111101010111011101000111010001010111010000011101000011011100001111000000010111000101111111110000010100011111000111,512'b00110001110000000111010100000001001111000101000100000011000101110101001111000000110000110100000001011100010000000100111101000100010111011100001111110101111111001100000100111100000101001111010001010100001100000100010000001100010011000111110001010100110101110111000000010011000101011100111101010001010100011101001101001100000000110000010100010001000001000001010011011101000111111111110000110111000000000101010001000011010011110011110001111100000000000100110101010011000100010001010011000000001111000100011111000000,512'b00000100110100111111000001010011000001111111010111000111010111000001110100000011000000010011110000010100110011000000110011110100001111011111111100010001110101001100011101110111010100110011001100010100110101000001110011111101110000001100000001111100110000010111111101110111000011010001011111010001010100000011010100110001000000000001010100000101000001000111010001111100010100000011000001110001110111000000010111010011011100110000010100010111000111000000011111000100010111010101000011000001010000000000110011010101,512'b00110111010100000001010011010011000001000101010011000101010000011101010011011100000000111100111101110111001100110100011100001111001111111111000011110101110001011100001111000001110001110000110100011100011111010100010100011111010101011101110001001111110000001100011111010000010000110001000111110101110101011100110001110001001101110101000000110100111111011101000011011100010100010011110000001111001111111111001101010111111101110000110100110000000111010011010100000000111101011100110101110111011100110011000011000011,512'b01010111000000000000000100000000010000000101010100001100010100011111000100001100010001001111000100000101001101001100001111110001110000000000011101000100011101110101000000000000000011000011011100011101110001000001010001000100000001011101111111011111001100000000000101000111110100110100000011001100110011111101110011011111110100000100000111110001010100001111010100000011000000010111001101011111000011011100000111001100011100000000010111010100111100110001010100011100001101110101010011011100010001110111010111000111,512'b11010000000100000000000001001111111100000001010000001111011101111100000000011111111101000101000101000111001100111111001101000101110111110100111101001101110100001101010000110100011100010001110100010001000001110001000101000011011101111100010111111111010111000000000001000000000001011101110000000000010101110100001100111100010000000000001101110100111111001100010011000111010000001101011100011101111111111111010111110000110000110111110011010111110111110000000000111101010100010101000100110011110001111100001101010001,512'b01010101110101110101110100001101110111111100010100010000000100110000000000000001111100110000111100110000111101000111000011111101010101000011000100110100111100000111000111011111110001000100010100000011001101011101000000010100111111000011110101110011000001010111111100010100110011010000000000000011111101000000110001011101110011011100000001010101000100001100110011000111110011111111010111000000000100011101111111110011110000010101010111110000000101000011110100000000111100111100111100111101011111110111111101011111,512'b00000100000011010100010011000111000111010111001100011101011100000111111100001100001101001101110111110111001100010011110101010100010100110001010100110100111100000001010100010000011111011100111111010100010101001101011111000100000011111111010101110000110001001101010001000001010000111100010100000000000011111101110111110101000011010111000000110001110011001100010100000100001101110011010011000011010100001100011101010000110100000011010111110101001111000111000100011111000100000100110001111101000101000111110100001100,512'b01000101010111001101000101110000000100011111111111010011000101001100111101000101111100110101000001000101010100000100010000001101010000000001000100010111110001000111110011011100000000001111111101011101001111001100111101110001110101111101010100011111110100110101111101110100000001110001000000110101110000011111000100011100000000111111000011001111000100010111000011001101110000111100010001110000110011110100110101001111110001010000110101001100110000010011111101011101010101011111110001110000110011000000110001010100,512'b11110011000101000101110100011111110000000011001101000111000011000011010001111101010000001100110011010111110000110011110011000111000101000011010100001100000011000111110100010000010000000000111101111100010001111100111101110000000001010001111101000011000101110111000101000000001101000100001100010100110011000111000100010100010101110001110000000011110100000000000111001101000000011100010111110111000000110111000111110101111101010111011101000100010001111101010000111101000001011101110001010011010011010000000011001100,512'b00000100111100111101111111110101011111000100010001010101000101110011001101000100010001010100111101000111111101010100000001010000110001010000110111011101001101001100011100011101001111000101000100000100000101011111010000000100000101010001010001010100110111110001000100000111110100000000110111010111000101110011111101011100000001110100010111000100110101011111011100011100011111110011011111000101010101110100010011110001000111110011000011010100111101110101110101110111010100011100110000110001000000000000000000010001,512'b01110011110000010001001101000111110000110011010001110001000100010000001101000101111100001101000001011100110101110101010111011100110100111100000100111100011101110000010011110011000011000011000111110011001100011111001101010100001100000011001101000100010100110100111101111111001101001111000101110101110001110000011111110100110000010011110111110001110011001100010111010011000011110100000000110011111101011111000100110001110000011100110011110000110100110000010000000001000000001100110000000101011111010000011100010011,512'b11110000000001110101110000010011010111110001110101010100000011010101110101001100001101000100110011010011010001000101000011011101110000011100111101010001011111010111001100000100001101001101010111000100010100001111000100000100010000110101000001010011110011010011001111010011010001011101110000110100001101010111111111011100010000110111111111110101001100110101000100010111010111001100001100000000111111001100000000110100010011000000001101111111000100110000000101110000001111111100110101110101010000001100000001000011,512'b11011111001101010000111101110011110101000111010001110001000001011111010001000101111100010101110111110111011100001100011100000011111100110000001111001101110100010011000000011100010000010001110000111100010100111100001101001100000011110001011101111111000111111100110001010000000100001100000111001100000001000001111100110101010111110011010100011101000100011111000101111101000111011100011100010100110101010101000001010000010000000001000001000100110011110001000100010001111100010111010001011111010101110001001100011100,512'b11111111011100010101000100110100010100000000000011110001000000110111111101010000010000000100110100010000000100010101000100110000110100110000111100110101000001110101111111000111111111010011000011110101010000110101000101010111010000001101011101011111000011000000110100011111010001001111111100001100000111000011011100000000110000010001010100011111110111010011110100000001000111110001000011110000000111000000010011000111111100110000010101010101110001000100010101000011010101000011010000010111000101000011000000110001,512'b01010100010011000101110000110111110101010001000011000101011101000100010001000001001101000100110001011100011101000111000001001100010100000111000100110000110111111111000001110000010011000011011111111111011111110100000000011100110001110111010011010011011111110000000101110001000000000101110101110011000101110001000100110111010100110001110011110101000011000100111111001111000011110001011111000000110100000011010111001100110001001101000111000011000101110001010001000111001111000011011111000101011100000001010101001101,512'b00000000010001001111010000110000010011000001110001110101000001111100110101000000000011001111110001010000000111001111000011110001110100110101111111110001011111110001000111010001110101000000001111010101110101011111110111010101000011111100000100010111000111000000001100110001000001111111110000011111000011000001000101000001000100000011010001011100110000001100111101110100000101110001010001110101110011010100110001110011000011010011110011110100000100000011000001011111010101000001110100011111110111111101110000110001,512'b11110000111100001100110000111101000011011100000000010101110111000101010100000001010100010001110011000111010111000100010001000000111111010001111101000001110100001101110101110000010111011111110001011100010011111100000000001100000100000111000011110101001111010011010101110111001100010001000100001100000000110000111100110111000011001101010000000101001111010000110111010011110111010101110100010000001111000101001111010111000101000001110101010101001100001100010111110111001100111100011111010000001100111100110011001100,512'b00001101001101010011110011110001011111010100110011111100010000110100000101110100010100010100010111111101110000001101011100010100001100010011000100000101110111110101011101010001110000111111010100110101110001001100000001000001011101110001010101000011110101110100010011011100011101000100000001010000110100000001001100110001110000010111000011111111011111000011011111011111010000000100000111011101000000010001111100011100010000110011110101010011001100110011110011110000010100110100110101011101011100010000010011000000,512'b11010000110000000011111101001100000100110000111111110101110101111100010011010100110100011100111111000000111111000111010100010111010101110011111111010111001111111101010011001111000001001100111100110011001101110001010101000100011111000000111100010111010101111101010001000001110100110100010011000111000001110000110100000000000001110011011100011111110100000111110011000100000000110100110000000111001111000011111100110011001101000011001101000000000111000001001111010101110111001111001100000111010000010001010001000011,512'b00011101000000000101001111110011010000000000111101010011001111000011110111000011000000111100110001001101000001110101011100110011010000010111010011001111010011110100010101000001000000010011110101110100011101000001110111001111110001011100010101001101011111001101000000001100110101000001001111000011001101110111010000000001000111011101000111010100110000011100010001011100000011110100011111010001010100111111110001110111010101000101111111111101000000001100001111000101000001010001000100010001010001010111111111010101,512'b11010101001100111111010000110001110100110111000111011100001111111111110100110011110000010101000000111101000100001101011100010101001111000011110001110000110001010101000011010000110100000000010011001100000000110000110011110100000011011100110100000011110001001100010100010100011101001101000011000000000000010101010100000111110101010001001101110101001100110000011100001100000100000001000011000000001111001100010001011101001100010001111100000101000011110011111100001100000000110101001101010000111100011100011101010001,512'b01001111000111110000001101000101010011000001011111000111000100000000010011001101110111000100111111001111111111000001001101110100000100000100110011111101001100000001011101001100011111000100010100011100010100011100111111000001111100000011011111011100010001000111010000010000011100111111010000111101001100110111000011001100001101000100001111111101110000010101000101000101110000111111000000010111000001001100111100010000011100110101000111001101000001111101110000001101011101001111011100110000110001000000110111010001,512'b01011100000001111101011111110000110011001101110111111100011101111100000001111100000011111100000100000001011100111111000001001100010011110101110000010000000111001111010101010011010111010100111101010001000101000100001111000100110001010101111101010011000011011100010001110001010111000100010000111100111101000011011100011111000100001101110001000101011101011101000111001111000011110000000111000111000100010000110101000101011100111101111100001101110000000000001101010011110001000001000100011101000000010100000001110001,512'b00111100010101010000110011001111011100000001000000010011111101000001111101010000000001001111111101000000000101110101001111011100111100010100000111000000110111111111000100111101010011111101110001111100000000110111110001011100010100010100001111010011000000000000001100010000111111110000010011000001010001000100001111111111011101010101110000110000001101111100110011110000000011111111011101001111001101111111110011110011010000000111110100010100001100010000010101000100000000010001000000000100110000000000111100000000,512'b11011111001101000001110111110111010101000001110101010111011111000000110100110011111100011111111111010011000101110001000111110011110000110000000101000001011100110000011100110001010011001101000111000001001111011100010001000000110000001111001111110001000001110001000100110011010000110001010011001101011111010011000100010011011101001101110000010111010100010100011101110001000100010100010011000001011101110000001111011100010101110000110001000111010101011111110000111111000011110100010101001111010000110101000100001101,512'b00110000000101010111010001010000011100011111010100001100011101011101010101110000001111110111000111110111010000010001011100000000110000001101010001001100110011001100010011110101110100010000111101010001000101000011110100001111000100111111110001110001000001000101110111001111011100000100000111110000010111000000110000001101011111010001000101111111011101011111000011000000111100001111010000011111110111000011001101111100000011000100000001010101010001001100011101001101010111110011110100000100001111010101000100001111,512'b01110100001101010101010000000000000111000011010100111100111111000101000011111100111100000011110000110011000100110111000001111111001101001100000001111111010011110001010100110001001111000111111100010101011100000001000000000100111111000111011100000100011101000100110001011100001111000100001100011111010111011111001101000101110000000000000100001101011111001100111101110001110111011111000001010101010000000000000000001101110101110001000001110101001100000011000111011101001111111111110111000000001101010001000000010100,512'b11110111010011110101010011111100000100000100110011111100000100000000001111011100000100110001110100110100010111110001001100110101110000110000000000111101000011011101110100000101110100111111000000010000110011000101011100011111110011110001011101110111110101001111111100110011000001001100000100001100000001110001011100001100010111000011000001010111011101000011001101111101000111111111000101010111010100010000000011001100000111110101000001010001110111000101000001010111011101111100110011010011110011000111000011010000,512'b00000000001100010101000101000101010001110100000101000100110111000011011100000100000011011101000000000100000000000000000001110111010000000001110001000000111111000000000101011101001111000101111111011100000100110000110100011111001100110001010000010111000000010011000100111100001100011111000101010001001111011111011101010001010100110101001101110100000011110111010001011100110011011101010000010111110011001111110111110011000001010100001100000101011111110111000101011101010101010111011100110100111100110111010111000001,512'b11110001111101111100110000010101110111000000111111011101000111001111000100000100110000011111000001001111010000010111000011010000110100011100010001110011000000010011010001000001010111000001110000001100000001010011000000111100110101001100010001001111000001110001010101110111010001010001010100000100110000011111110000110100000000001101010101010000110000110001011111010000110100110000110000001111010000111111110011010000011111001111011111110100001100001100000100010000110100110000010101000001010111010100111100111111,512'b01111101000011000001000100110011001100001100010001010000110011011111110001010111110000010001000111001100001111110111111100110101111111000100010101001100111100110001000000111101000000010101001111010011010001000101110101000001000000011101011100010001000111010100010000111111110011110001000001110001000100000011011111001101111100010001110001001101000100010000011100110100110011010100001111000100000111011101000000010011010000011101110001110111000000000111011111000000110000001111000111111101000111011101000011110000,512'b01111111000000010001110100000001001100110100001101010001011101110001010001000111001101000000000111000001011111010000110001000000001101011111000011010000000111010011110001000111111111010101111101010001001100111111001100110011010100110111001100111101011101111100110011110001000011110111000000010100010111110001110100110011110000001101111100011111010111110001000000010001011111001101010001010000010101110011110101010000000000000111110011001101001100110111110000111100001101110101010001110001010000011111110011010011,512'b01110001111100111100000011010000111101000011010001000100010011110011000011111101110011110001010000010101110100010000110001010000010011000000111100011100000000010111000100110100001101000000011101010000001100010011111100010101010011110101001100110001010100110100010100110111000111110001000100110100111101001100110000000100010000010000000000011100000011010011000111000000110011110001111111111100011111011100001100111100110000001101010000001100110100010000000001110100110100000111001101111101010001010111001111110100,512'b01110101111111000101001111000011000111001100001101000101110100010000000100011100010100110100010011110000111101000111000001110000001101010111010001010100110001111100110000011101000100011111000001011111010111011101000100110000010100110100000100111111110001001111111100000000001111110000010001000111110000000101011111010100110000001101111111110011011100110011001100111101001111110001000111001101111111110001111111011101000001110100011100110101010101000101110111010111010100000100110100000011011111110100011101010001,512'b01001111110100011101000001010000110000111100111100000001001111000001000000010011010000110001001111000111010111010011011111111101000000011100111100010111000000010100000000000011011101000001000001000011010000110001110000010011011101110001110101010101111111110101111101110000010100010111110100000100011100011101000001001100010001110011000011010001011111010011011111010101110000010100011101010001000111110100000000110100000101011100110111010001111101000101110011011101110000011100110000111111001111010101110001001101,512'b01000100010000010101000001010001001101000101000001010100111100111111000011001100010100010100011101000001000000110000011111011111111101110001011101110100110111001101110111000101000111110001110100010100000001000100000111010000001111000111000100000100110000110011110000010101110100010111010100010011010001010111110001011101001100000111010101000000000100010001110011010111011111011111110111010111110111110001000011011100010100000000110000001111011100010100111101001100110001010000000100011100000000111100000011001101,512'b11111100110011010001000100001101110000000111000011000100011111000011010100000100111111010000001111000100010000111100110000010000110101010011110111000100010111110101011101010001011101001111000001000000011100000011010100000101000101010011001100001101110000011111011111110101010111000011001101010000000000000100111100000101110000011100000000011100001101110111000000000001000100000011000000000000110001000111111100001101111111000000010100010101011111010011000111010100000011110001010011001100111111000001010001000100,512'b11001111001111111100000000001100110011110001000101011111000100000100111100000001000100010101110011000000110011111100110101111111010101000100111100010111000011111101110001011100111111000001111100111100010100110101000011110011110101000011000100000000110011000011010000011101011111000011010101110100110111010100110101010000001100000001010101110111011100011111110101110001010100011101001101001100011101010101110011110101000001011111110001000111010011011100110111000011000101001111001100110000000100110011000000001100,512'b11000001011101000101000000010111010001010000000100000111000011010111011100001111000001000111010001111100110100010100010000000000000101010111111101010101000011110100111100001111111101110100011101010000111101001100110100001100110011001111001111011100110001110011000001111100010101000000010000001101010100000000000000010001011101110101110000110111001111010001010001110000111101000100001100110011111101010111010011000001111101010111110001110011010100000000111101000001010100000011000101010000011100110100011111110000,512'b01011101110100000001000101111101000000001101010100000101001100010001011101000111111100011100110100110101000101010001111100010001000001110001111101001111000111000000110111000001010101001111000001011100001111111100001111011100110001110000001111110000000001000101111111001100010101111100000000000011001100001101001111001101110111111100000101110011110011000000111100111100110111000011010111110000110001001101010101111100000101011111010000111111110000011101110001011101111101011100000000001111111100000111110000111101,512'b01001101000100010000000101000000000001000011010001111100010000010111110111001100000100010100010001010011010100011111000000110100001100010101111100110001000100110101010111010011110001010001010100011111111100000001011100001111000100010100001100110101111101010100110000010011111101000000110000110100001111010011000111000101111111000000010111010000111111010101010000110011110101011100111111010011011111110111001101000011111100001111110011000100001111110101011111010011011111000001001101000111110101111100001100000111,512'b01110011110000000100110100110101011101000011110101110000110001000100001100001101000111010011000001010001111100001100001111001111110000000101110100011101000100110001110111110111000111001111110011000000010011111100010011111100010011111100000000000111000111000001010000000111010001110001000101011111110011111101110001111101111101110000010001000111000011000101010011111101000011110011111100000100111111110001001101011111110111001101010000110111000000001100111100010011010111000001001111001100111100001100111111000111,512'b01110100011100001100001100000011010101110000010100000001010101111100010100010111011100000011010101010101001100110100011101110001110100010000010001000100011101000011001100011101111100000101000001001100111111110011000000110000000101001100000000111111000001000101110100000000010011001100000000001100110111010001110101000000110101111101000100110100010100001100010011110011010111000111011111010011000100001101000001110111010011111101010100110011000111001100111111000101000000010001011100110011011111010100110100011111,512'b00010100000001010011000100111101001100111100110111010001001100011100001101010100111111110111110111110111000011110011000100111100000100000111010100001101000001000100000001000100000111111100110100001101011101111100000101010000110111001111001100010000001100000011011101001111110011010000111100010111001111000011000101010111110000000101110000011100110001010011110011001101010011010101000000000000010111010001110111110100010011000001110000110000011100000101010100110100000000011111010000010011111100110100000101110000,512'b00010001110111111111011100000000010000010101110111111111000101001111110011000011011101111101011101110011000011000101010101111101110111010001111111001111110101110111011111000111010000000101011100010000011100000011111101000011111111010101010100011100011101010001010111000000000000010000110100001100000001010111010000000011001100110100000001110100110000110000110011001100000111110011111101001101110011010001000001110011011111110011000101000101011111000000001100000001000001010000000100010000001101011111010101000100,512'b00011100000001010011111100110101000100000111001101000011011100110011011100010101001100010100010101010101110111000001111111010011010011110111110100000011110000010011010011001111000001000001010000000011000011001111000100010011000100010000000101010111010011011100111100011100000000011111010000000101110011000101010111000101110100010000000100001111110101010100000101111100011100001101001101111100000101000101110000110101001100000111010101010011000000110001011111110101010111001100000000110001001100000000000011000001,512'b01010100010011000011110001010100010101110001000000110100111100011100000000001111010000010011001101010000000001000011001101111101110000010100000100110001110001110101010011000111000011111100000011000111110000110000000000110000011101000101010000011100110100010001000011110011110100000001011101110001000100010111011101110011000011000001110011011111010111001100000011000001000000001111010111111100110011110011000001011100001101000011010100000011111100111100000111001101010000000111011101110000111111110011110111011101,512'b01001111010011110100000000000101111111000001011100110100000101001111011100110000110000000001000101001101111111010011000001111101110000111111001101001101010011010001111101000000010101110000010101000100000011010101010000111111010100110000111100011100000101001101111111010000000111110101011100000000001101000000011100010001110000000101110100110011000111010111110011010000000100000000000100000100110011000001010101111111110001111111000001110101111101010111111101110000001111010001000000000101110011001101010011001111,512'b00000000000111010001010000010011010000111101000011000011000001010000000100110111000001001100110100000000000100010001000000011111111111000101010001111101110011000000000100000001011101110011010111010101111101110011111100000011010001000101111101110000110001010111011101110100110101110011011101000111010101110001110000000000111100000111110111011100010101000100001100000011111101111101010001110001000001110111010000110011111101000111110000011111010100110000010111110000110111011101010011000100010111110100111100010101,512'b01010011001111010011111100000000000001010011000101010011010000110101000000011100110111000001010001000000110000001100011100000101001111000100010101000001010011010000110101010101001100010000010000011111110111001100011100011111011111011111010001000011110111110000010011111111010000110000110111010100010001001111010001001111011100111101001100000000000001000100001101001101010100011101001100001100000100011101000000000011010101011100110100111111000011110011110100001101110011001101110001111101110001011100011100110000,512'b01011100010111000100010001111101111100000100001100110001110100001111010011000100001111000100110000000000110011010101110000111111001101001100011100011101110100000000110100000000001100000011001101111111110011010111110000000101001101110001110100110000010000001100111100001100110011011111001111001111010011000100111111000000000100111100010100001111110000000011110111110001000100001100110100111100110000010000010001110011010100001100000011110000110100011100111100001111001101011101010101001101110111110111010011110100,512'b11010011000000000101010001000111110011011101011111110001010011010001011111000101110000011111010000000101001100001100110101000000000001010000001101110011110100110000000101001100001100000011111111011101011101010011110111111101000000000011001111111100000000010001000011001100011100111100011101111100001100010111000111011101000101110000011100000100111111111111111111111111000011010100011101110111110001110111001101001100000000001100010101110000000101010011110100001111110111110011110111011101110001011100110100000101,512'b00000000110000000001110100000011000011001101000001110000110001010000000000000100111100001101001111110111000101110001010001111100110101111100010111111101000000110100011101000011111100010011011111001100111111110011110001000000000111110111010100110011000111110101000100110100000100001100001101000011110001001111110100011100000000010001010101110001010011000000110111000011110011001100000011000001110101010000000100110011000101110000010000110001000001000101110011000001010001110111010011000111001101011100000111011100,512'b00110101010101111100001100000101000001010101011111111111001100000001011101001100111111000101110011110001010011000000000100010001000001110001110001110000010100000000000011010111001100001100011101000001001101000000110101011111110001010100110001010011010011010101010000010000000011110001011100000011110111110111010000001101110000010001000111000000001101110111111101011100010011000100011100001100001100010101010011000101110111111100010011110001010011111100000101010000001111001111010000010100110101000100000111000000,512'b00111111000111000001110001011101000111110100000001110100000001011101111101110111000011001100000101111100011100111100110001110001001111110000000001111111000111000011010111110000110001111111110001000001000000011100010000010100001100001101000011001101010001011101000000011100110101110011010101110100110011000000110000000001000000010111110000110100111101000000010000000001000011110111001100000000010000111111000000110000000001000011011100000101000100010000000011011100110000000101000011010011111101110111010000111100,512'b00010101110100000101110001000111000000001101110011010100010011000101110111111100000101010101000011010011010001000111001100000101011111010100001111000000110011011111010011111101010111111101010011110001010111111100110000111100010011000011011100010011001101010111000011110111001101111101000000110001110111111111110100011100000001011111000000010000010000110111010111110011001111000111001101110000110100000111000001010101000000111111110100010011000011110100011100110100011111011111110100111111111111110000010100011100,512'b01110101010111010101010001110011000011110100110000011100000011110111111101010001001100111111110100010011000000110000010011000101010011010111000101001111000100110001011101000011000111000101110100000111000001110011010111110000010100110101111100010001111111000000110001010100010111010001110001000000110101110001111111011100010100000001000101011101010100010101110111010100011100001101000001000101110011000000111100000000110111011111011111000100000001010000000100110000000101000000010000110011111100011100000111010100,512'b00110111110001110011001100111111000011001101000001110011001100000101110000000101011101000011010111001100010011110011000000001101111111110001001111000001000101011100000101110100000011000000001100000011010011011111000100011100010101001101000101010101110111000101110011111101111111000001000000000001110011001100000111000101110011001101001100010001010011000000001111111111110111010000000100110101110100011101000100000011000001001100010000011100000001001100000100011111001111001111000011110100111101010111011101110111,512'b11010111010011000111110011010101010100110001000011000100001100000100000011110001011101011100110111000100000100000111010100010011010011011100010011011101010111011111010000110100011101010101001111000111010101000001000011000101110000010111010001111111001101011100000001010001110001010011110100000001011100000111000000110001000100110001110100010011010000111101000100011100000111000000000011010100010001000001000000111101110100000111010000001111001111111101010000010111111100000011111100010101000000010001000000000001,512'b01001100111111110111000001011111000001000000000011011111000101111100000000111101000001000101000100110000000001000001001100111101000101010000000111000101001111010001000000110000111101001101000000010100010111000111110111000001001111010000011111000111111111011101111111001111000100000011001100010000001111110101110100110101011111010100010001001111000101000111011100001111010111000111011101010111110111111101010011011101001111000101000000010000110101010111010111010001000101000000011100110111000001001111001100010100,512'b01111111000000110000001111010101011111000000110100001101010101011111000001000100000000001100010001110001010001110001011101011111000000110000000100111100111111111100111100110001111101000101110100111100010100010101111100010000010001000101001100000100001100010000011111010011011111010111111111000011001111000001000100111101111100110011000000000000010001010000000000010101001101000001110111110100001100000111110001111111011100000100111101000111010000000000001100010000110000000101111100000011110101010011000100000000,512'b00000100011101000001011111001101111111111100110001000100010101110001000111110011010111111101010000001101001111111101010001001111111101111101011101011100000011111101011111001100001101110000111100011101010100000001000111000111000101001111000011010001010000001100011111000101010000010100010101000000011101011101010000111101010011010100000001110111110011001101011100010101000111110100110100001111111111001101010100000011001101001101111100110111010001000001110100000011110011000100000011000000000101011100010000000111,512'b11000000000011000100010100110011111100001111000000111111111100000100110001000111010100010111000100011111000001111101000011010011000000011100110100110001110100010100110001001111011100001101001100010000110000111100000011110001000101010101110011000101011100110000111101010000111100000011110000111111001111000100010101110000011111111101001101110011001111010000110011010111000101010000011100000000000000010001001100110101010111110000000111010001010100001111000100000011011111000001011111000000011100000000110000111111,512'b00000101010100000101000100111100010100110100000000001111000011110101011111000101011101000111110001000011000001000100000101001101001111000001011111110111011111010001110001111101000000110100001111011100110001110001000001110011000011010011110011010001000011110111110001001111110001010001000111000101001111000101010011110011110111000011010101000101111101110000010001011100010001010100110001110100111100010100000001111111111100110001011111000011001111000000111101001111110001111111000001000001000101000001110001010100,512'b00000100010000110000011100010100000000000111111100110101011100000100010011010001010000111100000001111101000100111111011111000011000111010000000000010100110011011101010101000100000101001111110000110111011100110111010001010011000101001101110001001101010111011101000000010000110100110011000000000011110101000001000011010001010011110000010101000000000011111100000111010001010000010101000001000000011101110101010100011100000101010001110000000101001111000000110001110101010011011101110000011111010001010111000100110000,512'b00010100110001110101110101111100110001000001110000110001010011110011011101110101110011111100011101001101001101010001000000110101000100010101011101010000110100110011000000010011001101011111000111000000110001001101000100000001010001001111010101111101110011010001011101000100001100110000010000001100001100000001001101000001011100000101111100010101010001001101000011001100111111110101111100111100110111001100001111110100000000110001010001110100000001110001001100111111111100111100110011000000011111110011110011000100,512'b11001100110000001111010000000001011111110011011100000101000011011100000101000101000100010001000001011100110011000001010011011101001111001111001111110000000001010001010101110000110001110111010001110111111101010011010000001101110011110011110001000000010101110011111100001100000011000000010111111100011101001101010101000111110000010000001100110011110100000011010101110100111100001101010000000001000101000001010001111100001101000011010001000001110000111111001100000101110100011100111100001100000100010000000101010001,512'b01001100011111000011110111000100001101010001000000000000010000010001010001000001010100110000110111110011111101010001000011010001001100111101011111010011011111001100011100110000110011010011011100000100110111011100110000110011111100110000110001000001001100111111000100010100111111011111000001001111111100001111111101001100010111110001001111010111010101000101110101000000010101010011000001010011000000000111001100010000111101110000010011000011011111010000010100000100110101010111011100001111000011000001001100001100,512'b11110100000000001101110011111111010111010011111100111101010100010100010011000000110000000000011111011101000100110000110100000000011111000011010001000000010011001100110101110011111100010100010100000001111111110000001111110011111101110011001111010100010011000000010001011111110000000000010011000000000011110001110100010011110100110101000000000111011100000001010111000101011101010011000011001111011111111101011111011101000001000001011111001111001101110101110100010001010101000011010100001101010011001101110000010111,512'b01000000000000000101010000110000111100010100010011001101010101110011001111001100110101110100000111000000011101110101000111010000000101010000000001110111000000011101010001000000011100110101010000000001111111111101111101000011010011010001111100001101111100001111000101010100110011011100010111001111011111110100010000110111111101010100000100010100110100110111000001110111000011000100010100001100110011110001110100001111110000000101011100010011010000110011010001000111000000011111010000110111010100001101110011000111,512'b00010101010001010101000001010101011101111100111111011111110000001111111101000100010100011101000100000011110101000001000001001111001101111111111101110100010111001111011100110001110100000011010101010111111101110001010111000011010101110101001101001100110111111100000000010000000100000100111111010111001100110001111100001101010100111100111111010101010111000001000111110011110101110011110100010001110000001100110000000000010100010111001100000100010100110100000100111101000001000111001101001100000101110100001111011101,512'b11010011000111000000001101111100000011111100010100011100000001010000110001000100110100110000001111010001010111001111010100110001110111111111110001110111001111111100010100010101001100000011010100001101000100111101110000000111011100000000011101000001000011001101010001010100010011001100000111110111110101111111000100000000010000110001111100110100000011000100001101110100000011000011000000010011001101010011000000010101110111010011111100010111011111010001111101000100110000010111000001011111000101000111010011000101,512'b01000101110001000100010011000001000111000001010000001111010011010111001101110000001100001100110100110100010000010111010100110101011100000101110001000111011101000101000100001111111111000011010000110001110000000000110101001101000101010101110100000111011101010101010001001111000000010100010111000001110101110000000001010100001111000111000111001101001101010101001111000111011111000101000011000000110000011111111101000001000000010000010011001100000000010100001100000001000100000111001101010000000011000001001111110011,512'b01111111111100011101010001001111110011010000000111000000000011000111011100010000000011111100110001010011010001010011001100110101010000000101011101010000000001000101111100000001111101000100000111000111110011010111000100111100110000110001010011000000111111110111001100110101110101010011001111111101011111110100000011110001110001010100010001000111110001001100011111001101010100010001110000111100011100000000000100011111000001000111001111001111010101110000010000000011010100010100000100011100000100000101000011001100,512'b01001101011111110001000001111100000001110000001100110100010100010100001100111100000001010011110100110001001111111111110000010001111111110001000001010001000001010001110000000011111101010111001100010011010001000000110011110011110100000001000011001100011100001111011101110011000000011111000001010000110101001100110100110111110101001100000001110011001111000100111111001100001100111101110001110000110111011111001111011100000000011101110101000111000011110000010011011101111100011100111111010001111111011100110011000111,512'b11010111010101001111111111110101000001001100111100111101010011000000011101110101110000010111010111110011010001001100110001011100010111000000010101010111000000111100000000011111001111010101000101110111001101011101001101000011000000111100110101111111010000000111110000011100000111001101010001110011111111010100110011001111001101111111000001010100010101000101110100011100111101010101010101000111111100010001110011000001110001000101110101011111000100000000010101000001001101010100000111000011110101111100010000010001,512'b00001101010000110000110000000100010000001101000101001101110000111100000001010011110101010101000100000011110000110001111100010100000100110111000001110111110000000000110101011101010011010000010011000100111101111101010100110100010011001111110111000001000011010101000001110111001111011101011101110000110001000000010101001111010000000000110111010011111100110111000100110001010001110100000001010100110000001100000001010000010100000111111100000100011111110011010100110101110000000001010001010101000011001100111111000000,512'b00001111011101000111000001110011110111110101000001000011001100110000111100110001010011000001001101010111111100010001010001111101110101010111001100000001110000000100010011111100110001110011011100111111000100000000000100011100010111110111001101000011010001110101001111110001110101010011000111001101111101110011110111110000111101000101000011110111010101001100001100110111110001001111010011001111111100111101001101001101010001000100001100110000000001111100001100110100010011010011110011010001010111111111000111111101,512'b00111111110100110111010000001111110111001100111100110001000001110011000001000011000100110100001100000000010000000001000001000001000011000101111100111111000001010000010100000001001100110011000000001100001101110101110100110111111101000000011101110011010000111100011101010100001100110001000100010100110001111100001101110100110101000000000011010000001100110011010001001100000000001101001111001111000111111100111100010111110100111111110011010001010100011100111111010001110101000011001100010000000001110111001111000101,512'b00010111010011010111110100110011000101000101110000000000010100010100111100000000110111110101000101000111110011000111110101010100000100000101001100001101000000010101000111111111110111010111010011110100011101000000011101011101011100010001011100010111010100110011000000000001010111011100010000010101110001110111010011010000010111000000111100001111000001110100110101001100001100000011011101000101110100011111110100010001001111000001000100001100000100111100000101110111001101000001111101010001000011010001011111001111,512'b11000000000001110000110001010001011100110011000011010011010100001101010000010100111101001101000111000100111100010011010111111101110011110001001101000111001100000000111101010000010011110111110101000000000011110011000000010001000001000001111101000000000001001111011101000001000000010101001100110101000000010001110100001100000000001100011101110011001101111100110111010101010011000111001101010000000111111101011101001111000101000000010100010111000101011100000111010000111111001101000001000011000011010011000000010100,512'b11010100110001000111010000000011010100000001011100000100001111010111000000010101001111000000111101110101000001000001001111011100000000000011001111001100110101001100000001011111001101010111010000000011111111001101010000000011001101110111110011110111010100110111010011110000111101111100111101110100000000011100111111011111000101010111000001010100001111011101000100011111111100000111011111000100000100010000010001000001000011001111111111010100110111010101001101110011000001000101001111011111000001110111010100000011,512'b00111111111111000101000101111101010111000000110001011111110011010111110100010100010000110111110001000101010011110000000000000100000100000111110000110000011101000001000000010101010111110001001111011100110011010111001100001101010000110101110001110100010101000101000100011111010100001100010000000000111111000111011101010000001111000111110000000100110111110111110011000011110001000001000011110111000011010101000101000001110011000000010101000111011100000101110111000001010000001100010001010111000111110100110000011111,512'b01111100010011001100000111001111110100011100111101010100000001000001010000110011110001110011110001010011001111111111000101011111000000001111011101110100110000000001011101000011000111000100000101110101110100011111000100000001000100010011111101000100010000010101110100001101110000011100010111110101011101110000111100011101011100000100000111010001110100110000110000000100001100000111111101110111111101010000000001010100010100111111010011110001001101111111000100000111000001010000110011010101000011000111000000001111,512'b01001111010101110011110111001101001100010100110111000101000001011101110000110101000011010000001100110101111111110011111101110000000001010111000111000111110100110101010011001111110100011101010100110100001111010101001100111101011100111111010101010100110101000001001101000011010001001100111101110011010001110100011101000000000101110100110101011101001100000001000001000111111101011100001100110001111100010000001100111101111111011101010000001101000100111101000001000100110111000111010001000000111101001101110111000101,512'b01011101000111011111110111010000011111001100001101110000110000010100000101000001000011000111010100011111000111111101010001001100110001001100010001001111010000111101110101111111110100010111001111001100110100110000000001111100010011011111000011010011011100110001110001000011000000110001011101010100011101011101110011110101010111111111010001011100010001001101011101001100011100001111001111110000110111010011011100111100111100110000011111111100001111111100010000010001110011110001011111111111111101111100000001000000,512'b11111101110000110100110001000001000100000011110011011101000111000011001101010000000000110000110000110100000100010101110100111101011101000111001101010011001111011101110111001100000111010100000000001100111111010111010000001101011111000001010111011100110001110100111100000000011100011100000001011111000001000000010000011101000000111111010100010001111100000100110001110000111100110000010100111100010111000011001100000111110100110011010111111100000100111100010101001111001101111101001111010000010111110001110100011101,512'b11110100000111110100111111111101001100000000001101010101110000011111111100000011110100000101111101010111000000000101001100000000000011010100010000110000000101111111110011000111110000010111001101010001110001010101011101010100010101000000010001111100000111010001010000001101110001001100000111110101110100011100000001001101110001111111110100110000001101110101110100110001000101110000000111010011010000110111110100011111001111010000110000110100000011000111011100000101110011111100110111000101110000000001011111010100,512'b11000101000100110101111100001111110000000111011111001100010111110000110100110011110000110000010011001111000000011100000100000111000000010111000000001100010001010001000101000101000001111111010000001101110100110100001111011101000001000100000011010011110000010001110011000000000100110100000000001111110101110111001101000011110001000011000001111100110011111100110100001100010000010101110101000011010101000000111111110111110100000101001100010100111100110000111101110101000111000001011111010101110000010111110101010111,512'b00111101010011110001000011010100110000011100110111010100001100010000000011010000111111011101000100001101111100110001110000110001001111001100000111001111000100010101000000010000011111000101000000010101111100011111111100001100110100010000010011001100000101000001001101110001001100010101001111000000000111010011010000110001001111110111110000001101000000110001011101000101111101011101000011000111010000001100000001010000010101001101110101000100000100000101111111110011001100111100000100011111110111010000110001000000,512'b11111100001101110001000101000101001111011111000100001101111111010001010001011111011101111100011101110001110101001100000011000011010001110111001111010011001111000111011111011111110100000011010100010100000001010100000101000000011100110100010001000101010001000011010001011101010111001100001100111101010001000111011101111111111101111100111111111111010101010101000100000011011101010111000011010000000011111100010001011101000000011111011100010011011111000000110001111101001101111100011111111101110111010011000011001100,512'b11010011110000010111000111010001111101011101010100010111001100010011000101010100011100011100000001000001001100000011010100000100000111000000110100010100000100111100000001000011110101010101000100000011001101011111000000110011000111111111010000000000010000000001000000000000001100000011000100110001111111001101000101011111000000110000010011110000000001110100000100110111000011010101010011011111111101111111000101010101010000001101010011110000000001000101000000000111011111111100011101111111111100010100010100011100,512'b11010011111101111111010100000000111111000000000100010000010000110011001100000011110100110011010011010000010001011111110100000011000001010011000001001111010001110001010001110000011100010011010001110001011100010001000011110011110111000000011100110011001100000011001101001100110101000101000000110001011101000100110100010100110011001101000011010101011101011101000000000111110011110001001111111100010001110101011111001111000001001100110111010000000100010100011111111111010011110001011111010000001100000111001111001100,512'b01001111110011001100001111000101110011010111111101010011000011110000010011000000011100111100001101010001000101111101000000010111011100110000000101001111110100000011000000110000110001000111111101000011010000010100001111010011001101010011001101110001111101010001110011011100110000000000010011000000110000110111010011011101011111111100000000011100010000000100010001110100110111000000001111010100001111000001001111010000111100010111111111110111000000110000010100110100110000000000110000000001000100000000010000011101,512'b11000001000001110111110100000001000011110100001111111100010000110101110011110000001111001100110100000111000011110011110000111101110011010111010101000111011111011100110000011100000000010101000100111101111101010111110000110101001111001101000000010001000100010111111101110111000001010100110001010001111111110111111101110011010011111101110001010100000011110100010000000100110001001111110101010011111111010000010111000100111100010011001111001101010001111111011101110111010001000111000000001101000000110101000000110101,512'b00010000001100000000010011111101011111010011000101011101111101110100000111001111000001000100111100010100011100000101111100000001010111000011000100000001000100011100111101111101010100000000111101011101010100010000010100111100001100110111000011110000011111010000000001000000111101110001010001000011110101111111010100000100111101000011011101000000000101000001000100010011001111000101000001001100000111111100111101110001110000110011001111000000000111000011111100000011110000000100011100000000110100011100011101110001,512'b00010001110000011100000111010100000011010111010011110111000100110011010111111100010101010001000000000001010011110011001101110111110001011100000100110001011111000101011111010001000101110111011100010101110001011101010011110000110011000000110101000011001101110011010111000101001111001100010101010011110000001101110001010111111100111111000001001100111111110111001111010101110100010100000001001101000111111111110100110100001100110101001101000011000011000000110001110001000101110001110011011111010100110111010011011100,512'b01000100110001001111000001010100000001010101110000110001001100110001111100001100011100110000110001000000111101000011110111001101000000010001011100110011010111000111110000000000011101110000110111110100000101000011000100010111001101000001000011110011000100000111010101110001011111001111000001001111110001011111001111011111110011010100111100110111010100111100110111000101000011111111110011111111110111110111000000110001110101111101110101010111110011110011010000000001010001111100010000010000011100000100011111110100,512'b01010001000100010011000111110100110000111100110000000011011100000011010001010000001101000111110101110011000000110100111100010011010000000000000101001100110101111100010100010100110000000000010111010111010011011100111101000111000011011101110011110001000011110011000100011101011100110101001100011100110101000001001101110000001101010100001111000100110001110111001101110001110100111111110000110011111101010111000001110101000001010101110100010000000101011101001100010100011100111111000101110101010111111100000111010011,512'b00000101110000001100110111001111000101110011110111010011000000000001011100010000001111110001010101001101001100000100111111111111111101011100010000000111000100000000110011010111010111110000110001000000000100010000000011000011010101000100110001110111010100001100000001110101010100010000000100010100010011111101010100000000011101011101110000000011010001010001000000010011000100110100111100111101111100000101011111010000001101110100111100110100001101000111010001001101011100000100010001000111001100010111111111000100,512'b00110101010100001111000111000001011101110011000000010000111100110011010000000001000101011100110011111101011111010000001100001111110101000100110101010011000001000011110000000100010011000000110111000100110001000011011101000101111111001100001101000011010111110111110101000001010011011101000111001100110000000001001111111101110100010111000101110111011101000000000101110001111101110101000000000100000001110111001100011101010001110011110000001111110111111111110101001111010000110001110001000101110000010100000000000101,512'b01010001011100010000000011000001000011110000000000011111001111000000111111110111010000000101000100010001000101000000110011010001110100110000110101010001110000010100001111110011001100110001000101000011010001110100110000111111011111001100010011000011110001111100000100010111000000000001110100010011001100000011110100001100000101111111001101000111010100111101011101000001111100010001110001111101011111010000110101110000011111001101111101001100010101001111111101001100011100001101011100110001011101000000010011110011,512'b11000111110001110011110001000011000000011101001111010000001111000101001101000000111101000011010000010011110000110011110011000000010100010000110111010111110100001101000011010001010101000101010100001101110000001111000100110111111111010101110000110000000000110001110001011100010001000001000001011101000001001101000001010000001100010001000000010011110011000100000100001100110001010001010000000000110001010011110000010100011100010101011101000100001100111100000000000111110101000111010000000011010001011111000111010111,512'b01010001000101010101001101110001010001111100000011110000110111110100110000010111110100011111001111000011010001110111110101000111010011110011001100010100000100011101110001010101001101001111110100001101011101011100111100010001000000000000010100001100000011011111111111110101001100001100110100001111011101000101000000110000010101001101001111110000011101010111001111010111000100010101010101000111010000110011111101110011111101010000010000001111000000001100000000111101000000110001110001111100111111111101000001110000,512'b01010011010011110001001100111101010100010001010100110011011101110011110101110000010000011101110001110111110111000011111101001101110001000001000101000111110101000001001101110011110101110011010001110100111100000111011100010000010000000011111101001101111100010101110101110001111111010001110001010001111100110100110000010000001101011100010011010000010100000111000000111100111101000000110111000101111100111101000100110100001101000000111100010100011101010100110001010100000001000101010101001100000101011101011100000011,512'b11000100000111000000111101010101000111111111001101110001110101110111110000000100111100111101110000000011110111110111010111110111000001000001000000000000000100000111001101011101000111000100000001110011010001110001001111010001001101110100010111110001000101010011010101010011000001110011010000010011010000000111110100110100001101010011011111000000000100110000000101011111111101010011011111001100001101000001000000011101000011011101111100010001110000001100000011001100110000000100010100110001011111000011000000000000,512'b11011101010001010100000000000000110011000000010000000101111101111111011100010000000011001101110111000001000111001101001111001111110111010101000000110001010100001100001111010001110001010000000000011111000011001100011111001101011100010100111100010000010001001101010111000100011111000011010001010101010001111101110000000111000100110001010000111101001101010000000001110101010000000111000000110001110101000111110101110100110000001111010101110000000001000000110101111100110001001100001101000001000000000100011101010001,512'b00001100000100001100011111011100000000001100000100010011011101001100000101000011010000001111110100001111000001111101011100110001111111001111110100010011110100000101110101000000111100010100000111110101010011010100000000010001010001000011011111111101000001110000010000110100000000011100010100110101010001000001010000010011110001111111011111110100110000001111010001110011010011110011001101111111000000110000111111000100010100000100001100110000010100000000010001010100000100010100110000111101000000000011111111110011,512'b11110100011100000001000111010001110111000100000001110100001101010000110101001101000111011100110100000101000101001100000000111111011101001100110100010000000100001101110111001101010001010001000001110000000100010100000011001101010011001100110100001111110011001101110011011100110001110101000011000101010001000011110100000011110001110100110011110011000111010011000000010100000001110000110100011111010001110111010000010000111101010011000100000011110001000111010000110101010111000000010000010100001100111100111101011100,512'b11000101000100000001000100011101001101111101110100000100011111000011000000000000110011010000011100010001010011000000010000010101010100010100001111000111010000001111010000110100001100110011111101000011010011111111010111000001111111000001000101000111110100011100000111001101110100000000000000001100010011010111110001001101000011001101110100111111010100110001000100010000000000000101011111000111010100011100111100010100010101010101010000111100010100110000111101011100110011000101000000011111110001111101010011000100,512'b11111111010101010100000011111100110101010011110011000001010011010111000001110000111100000001001100111111001100001111000001110011000100010000010000000000001100001101000111010001000101011101000011001100010111001111001101001111011111110001001101000000011111001100000011000011110001001100010001010100111100111100000011110100000001110100000011000011000011111100000100110000001111111100110000000001110101111100110001010000010000010100000000110100110111000000001111000011000111011111110101111111010011000100110111001100,512'b01010111111111010111010000000001111100110000000001010100010000010111111111110000011101000111110000010011111111110100110100001101000111110011010101011101010101000011110001000001010000110101010011111101110000000100010011010000111101001111000011000000111100000011000011000111000000010011011100000001000011000100010001010000000111011111001100001111001101000111000000110001110100010101011101010101111100010011110001010100110101000100000001010100001100110001110001000001001101111100000100010111011100010011010001010011,512'b00000011110011000011000001110101110000000100011101110101011100000001110011000001010000110001110011010011110000110001000111111100000001000001000101010100110011111100010111110100110101111111110001000111000100110011000111110001010011000000010001001100010001010001000001000000000001110011110011011101010100001111001100110100111111001100010100110000010101000000000101011111000111011111000100110000001101110000010000110111011101000101110111011100111101110101000000001111000001110000110111010100011111000011111101000000,512'b00111101011100001101010001001101111100000101000000010001000011110011110000110011111100000011011111010001001100111100000111110011000001110000110011001101010011110011110011010100000011110111111111111100111111010000111111010101011111001100110100011100110111110100010101010100001111001111000011010000000000110011010111000001011111001111001100000111010100001111111101000001110100000000000111000000011101000001110011000001111101011100111101011100011101011111000100000111110111110011111111001100111101000100000001000000,512'b00111100010000111100000000001111110101001111001101111111010111000101111111111101010000111111001100000111110000000000010011010101000011011111010011111101000001010011110011110100010111110001000001011111110000110111010101110111011111011101110111010100010111110001010001011111110101000101010000111100001100000000010111001101111101010011110000010001010011110011010011000011111111001111001100110000001101010001011101010000111111110011111111000011010100000101110001001101010111011111010000011100001100000011011101110000,512'b01001100110011110000000101110100110001011111001101110000000101000100000001111111010100011111001101000100001101110111010100010011010001000100000100001111011100010001010011001100011100110101011100110111110001000111010001110100010001011111110111111101000000000001011101000000010100111101010100011100000011110001001111000101000000111100111111010001001100010000110001000000110011000111010101010001010101010011000100010111001100011101001101000100110000010011110100010011011111110011110001110011000100010101000000001100,512'b00000101001101010111011111110011010101001111010000001100111101011111000111110011010100000101001100000100000001000000110101111101010111000101010011010101001100111101111101000011000101011100010000110011000001000101110011010101010001111101000001010001010000111111001100010100110000000100110011010000010011011100110101111111010000000011001101010000111100010111010100001100110101010000001100110100011100001100001101000011110100001111010101010111000111011100010111011111010111011100001101111100010000010001010101010100,512'b00011111000011110101110101000000110011000111011111110000110001001101001100001100110111011111001101000011110111111100010111001111010001011111110100110000000101000011010000000000110011011100010001001111000111000100000000001101011111110000110001010100000001010011011100000001111101000100000011010001110111000000011101110111110011000101010101110111001100111111000001111100011111110100010100110100000111000000000011010011111101110011001111000001010011010011110011110001010111010101000100111111110001001111001101010001,512'b01110011111100000000000000000011000000000011010101010100000111000000110101111101000000110000010101110001000001010111001101010100000001111100010101111111111101000100111111001111000100001100000001010000010111110001011111001100110100110101111111110000001111000111000111010011000000010011001111111101110101111100011100010011010111010100011111000101110001000100000001000100010000110011110111010101110000010111110100000000010100110011111101110001110100011100010100111100000100111100110111010111110011110000000000000011,512'b00110011110100110000010000110000001100010001110001001100000101110111000100001111000011110011110000000011111101000001000011000100110111000111010111000101000011110011111100110100110001001101000111011101010001001111110011010001000000000011010001010100011101001100111100110000000001010000000111000101010111000100001101110111111101000000000100010111000011110000000100010111000001001111111111110100010011000001000000110100010001010001011111000000111101011100110011110100010111011100111111010100001100001100000101011111,512'b01110000000001000111010001110100111111000101110101111100111111000100111101000001000000000111010011000101111111000011000000001111110001110101110011111101010100000111110011110011110000001100111101111101111111000001011100011111111101110000110011001101110101110011000101000100110111010001000100111100011101000101001100011111000011000001001100110000011111111111001101111100000100011100110001001100000011010111110100110001010100000000110101000011000100111100110100010101110011110101110111001100000111000001000001110000,512'b01011101000001110101001101001111010100000000010101000111010000010011000101000101011111000100011101111111110011000000010000001100111101011101000100000001000000111100000000000001010001110100111111011111110100000111000000110111111111010011111100011100111100000001010100010000000001000100000000110101110000010111010100000101110100110000011111000111110001010011110101000111010100011101010111000001110001000000000100011101111101001111001100110100111101010111000111010011110101111100011101110011010000110011110011011100,512'b11110000001100011101000011010111111101111101110101000011010011110001110100111100000001110000011100000111010111010100110000111111001111110111110111111101000101010100000011000111110100010111111100011100110000001101010001110111110000000000011101011100110111000011111111000111110111110001110001010100010111111100000100000000000101010001010100110101001101111100010011110111010100000000000001000001000011010011000000111100000101001101000111000000111101010001000100000000010001000000110001000001000100110001010100011100,512'b00000000110101000111000001000000010001000001010100001111000011001101000101011101001111011111001100011100011100010000010100000001001101000001010101110001011100010000010100011100111100010111000000110100110011010001110001110001000111001101001100000111011101111100010111110011000111110101111111011111000101000000110100110101010011011111111101110001010111110011010001010000010100011100000000010000001100111100111100000011111111110001110000110000001101000011010100000011000111110011001111010001010011010111111101001111,512'b01110000001101111100000100011111010001011100000100010011110100011111010000010001110101000111010101110101110111110000001100110011001100010101000000011100001100110011001100010100001101001101110101110000010000111101010101010000110000000100010011000011001111000100110001011111000101001100110001110100110111000111000111010001001111010001010011000100001100000001001111011100010000110011010100000101110000110001000001001100000011000111001101110101110011000011000111110101010100010101001111010001000000010101010001010011,512'b01001101001100010011010111010101001111000000010000001100111100110000000000000111010100001111000100110011000011001100001100010100110001000100010001111111110101010001000000001111010011001111000011010100010100111111011111001111001101110011110101001111010001010101000011000001000011110000010000010001000011000100111100111100011101001100001100110000110000000000000001000000000000010011110000111111010000000100001101111100011100001111110011110001010000111100111101000000000000110000001100111101110001110101110001110101,512'b11000000001100000001000100000111001100001101010100111101110011110101010101000100000000000011010011110011000000001111000111011111110100011100011111010000110101110001011111010100110100010011110000000100111101010111001101001101110000111101000111000111110100000100110000010011000011111111110011000000010000010000000100000000011101010111000100110101010011000000000101010011000101000100001101010100111101010100111111110000011111011100010100111101110011010011001101010111111100111100111100000111110011010000010101110011,512'b11000111000011010101000001000001001111010111000011001111000000000000111100000101011101110000001111011101011100010011111101010011001100001101111101110100000001001100010111010111001101001100000111110011001111000011010101011100010011111101110001000111111101000100000000010100001100010101111100000001110111011111010101010111010101111111000011011101010100110000010111110001000111011100110100110101010100000100110100000100010000011100000000000000001111001111011101111111001100110101011101000100010100000001010101010100,512'b01010001011100111100110001111111110111110100000000000011111100000000111111011111011100010011110111010101111100000000000000011101111111001101011111010101010101011101110011010111111100110011010001110011000100001100010111000100110101111100110101110111010001110100110000011100000011010111110100010001111100110011110011110100111100010000000101111100010011000011110101010101110100000111111100010111010011000100000101110100010101011101110011001101110000011111011101001101000100011111010100110011110111001111010011010100,512'b01111101110001110100000100011111000000110001011111010101110011110001111111110111001100000011011111110000010111000111111111001100001101110101110111011101010000011101001100011101000101111101110000000101110001000001110111001101110100111101010000011100001101000101001101000111000001000011110111000000000111000001110001000100111100000001011111110000000000010101001100000011010000110011111100111100000011110001110101010011000101001100000000011111010100110111110111110101011111011100001100110001110000111100000011010001,512'b00011100010000010011001111010101110000000000000100000001111100111111010011000100111100000001001101000101000011111101110000001111110111111100000001010011110000001101001100001101010011110000001101001101011111000000011101001111110011000111000111110001010111011100110001001100011101000011010100110100110011110100001100000001010000001111010101010001110011000100110100111111000011010101110111001101000111011101111111000011001101011111011100110000001100000111010001000100000111000100010001110101000101010001010101000100,512'b11001111000111011100010111110001010011110111000011010011111100010111110011000100110101001100111101110000110000001101000101110100110011000001001100001100010101011111001100000001111101000011001111110100010000111100000111000000111101010000000000010000000000000111001111010111011101010011111101000000110111000100010111000100111111001111000000111100000001010001010111110011000011010100011111110100001101000100000001000111010000010100000100010101001100110111111100111111110111011111010101011111001100011101011100111100,512'b00000011111100110000111100000111011111110111010100110011111100001101111100000001110101000100111101110011110101011100000100010100001111000100010000011111110111111111001111110101010111000000110001000100000011000111110000000001110111000001000111110000110111110000010011010011000011110100000011001111000111000100011101110111000111110001111101010101000100110101010000000011110011000101010001000111010101000100000100000011110000000000000001010100111100110011001111000011000100001101110101110001000000110101011111001101,512'b01111100001100010101000011111111110100001101110001111111010111110100011101001100000001000011001100011111000100000111000101000001000000010000000101001101010100000100111100000011010111000011110011001100010001010011000111010001110100110001110000010011010100010011110001001101000000011101001100110100011101000100011101111101111101000101000101110000010111000011011100001100011100010100000101001111000101001111010100000000010000111100000001000100110011110100000111000100111111111101010000110101111111111100010000001101,512'b01000100001111000101110100001101000000000001011100010101000000010000000000110001001111000111011101110101111100001111011100010100010000010101000000010111000111000100001111010100000100110000010011110100001101000101010111011100011111111111010001011111110101111100010000000000010011001100110100111111110011000111000000001111110000000011000101010000000011000111000111011111001111011101111101010100001101001100110000000011011101001100010111011101011101000100110001000111011101000011110000110011010111011111110101001100,512'b00110000110111000011000001110011110000000100000000000000010011000011010011111111000000000101110001010111000001000100001111010000110100010000000000000001011100000100000000110101111111010011110100000000000000110101111111010101110101000100011101001101111100000101010111000000011100110111110000011100011100000100000100010101010000001100000111001111000100010101000101000000110000001101110101110001000000010100110001010100011101000000000111000111111100000111111100000011110011000001110011011100000101000011000000111100,512'b01010001001101110011110001001100011101111100001100000011001100000000001100110000110111010001010000010000010011001100111100111111110011001100000111111100000100111100010100111111000000110001111111010011000011011101000100000111000000000100110000110111110000111111001101111111110101010011110101110101000011000101000111000000000101000001000000110100011100111100010100000111110111010001000101110001000000010101111111001111110100010111110100010100000001110000110100000000000001010100000001011100110111111111110101000001,512'b01000001010001110000110011010000011101011100011111111111000101000011000100001100000101000000001101110000110000010001110100110000110001010100010101000011001100000011000000000101111101001111010111001101000001000000000111000111001111110100000000001101110100011111000001000011000111001101000000001111000100010111110001110111010001001111010100010000110111110000000111001101000111110101110000010100011101010101001100110101000101110011000001000000010111110100110111001111110100000100011100010001000001010000111100010111,512'b11111100001101000011001100000000110011110111010011000101000111110101110000000000000000110000010001110111111100000111011100110101111101110100110011000001000000111101010111010101011100110100010100000000110001011111010100010111001111110111011101000000010000110001111111000101000100010000111101011111001100000100110111010111000100000111010100000100000101001101011100010011110000010011000111001100011111110111000001010001000100001111001111000011000000110001011100110011010001010000010011010000010111001100111101010000,512'b01010111110001000100110111000011010000110111010001011100110001001101110101010011011100110111110001010100000000001111000100110100110001000011001100110000000001010101000100001100000000110100110111010111000011001101001111001100000100001111111101000100000001110101001100001111001100010101111100000101111101000011010101110111010101011111010100001111000100010100000111010111010101010000000101000100010111010111111111010000010100110101111111000111110000000000000111001101110001111100000100010000000000000100010000000100,512'b11110101110101001100010101000001110111010011011111010101110111110001000100000100000101000011110111001100110011001101000101000111010001000100011101111111000000110001000101000101110111000111110001000100001100000000110001011100110001111100011101110011000000110001001100001101010100010101010000110011000101000001010000000101011100110000000101000101000101000001111100010011000000111101010100010000010001010111110111001111010011111100110100011101001111000100110000000011010100111100011101110111001100111101010000010011,512'b00001111011101011100011100010001010101000001000111010101000011110100000111011101111100110111010000000001110100000100000011011111000100010011000001110100000100110000001111011100000001000011111101000011000001000000010001010001000011000011110001000101010111001111010100000011001100001100010101110000110000010111110011011101010111011100010111010000010011001111000100001100000011110101001101000000111101111111110101111111001100000011111100000101000100000000110100111111110001110100000100011111110101111101110011010111,512'b01010100001101000000000000001101001111000011001111110011110101011101001100000111010000011100001100110100011111000100010001010011110001000100110101000111111100000111111111000011011100000011010000001101110111001100000011010100010000010100110111000001110101010001000000110000110011110100010001011100000111000100110001000100001111011100110000011111000100110111010111010111010100000101010011001101110001000000111111000101110100011101010101111100011101010101110011111101001111000111010011000000001101000000011111111100,512'b01000111010100000001010101010001111100001100011101110100000101111101011101001111010001010100011100001101011100001101010000010101110111110101010100011111011101000101010001001100000000011111000000110001001101110011000111110101110001010000011101010011000111110101000101001111000000000101110100010111110101001111110001110011010100111100001111111100010100001101110001000000011111000001010011000100110000010011000000010011001100111101000011010101110111110000010111110000111101000001010101111111111101010100110111010000,512'b00110001010000010000010000001111001101000000010100011101111111001101110101110011001111110000000101011100011100001101010101010001111100110100000111000100110011000000010111110100110011001111000000110100110001110100110000110111000100010111001111110101010000111100010111001111111100000011111100000100000100000100111100011101000111001101110111001101110000000001010111110111110001110100000000000011000011010101000111011111110000000011001111001111110001000001011111110100110101110001010100000011111100011101000000111111,512'b11001101000111000001000001001101000001110101011100000000110001111101000111000100001101000000001100111100001100011100010000000000001100010000011101110100110111110000001100111111000101010000001111110100011100010011110000000101010000111111010100000011110001010000000101000001000100111100110100110100010001110011010100000011000101110000111100001101000001010000111100010111000000000000001111110001000001010001000000110000001100010000111100010111000000011100000000011111000011110001000111001101001100000001001101001101,512'b11001100011111000101010000110000111100110001110011001111111101110111010111111101110101111101011100110111000100000001010011110111110111010100001111110000000111111101110001110000001111110111000101010001111100011101110001000111110101110101010111001100010000010101000000010000011100110000001101000000010011000001000011011101000011000101110000010101110100001111111100110100000101111100110000010000000101110000110001110001110101110000000000110001110001000001111101110001001111011100110011111111110100110100110000110101,512'b01010100001101010011001100001100000001110001010001000101000011110101000001000100000100010000010011010000010000001111111100000001110101010000111111110100000000000100010100111101001111110000000001001101000101010011001101010011111111110011010000111111001100111101111100010000010000110001001100000101010011110100010100110011000011000100110000111101010000111111110101010100011100000111000011110001000100000001000001000000001111001100010100000111010000000001010111001111110101010001000100001101000011011101000100110001,512'b00000111001101010001010100000001000000000100110100010011010011000100110011111111000101010000111111111111001111000001001111111100001111110011010011000100001100111111010100001111111111000000110100000111110001000011010011010111110111010111010001001100010001011101001111110111011100010011011111011111010101011100110111011101110000011111010001010100110101001101000100001100010011110011111101110100000000110000000111001101110100011111111111110011111100111101001100000100001100000011010101001111001111000001000111110011,512'b11110100110001001101000100000011110011000111010000000000010000000000001100001100000100111111010011000011110111010011010001011111010100010000111111001111000111000001000101001100110011000111010011011100010100010000110011010111000011000111000011000111000011000011010100010011000000110000010000110011001101010101000000011100000101011100001100010100001101110000000011010000110011000111111100111111000011110011000000000101000001010001000101001101010111001111001101011100011100110011000100010101110001111111111100011100,512'b01110100111101011111000000111100111101000101110000000001010101000101000100000011110001000111000111110100011100000001001101110000000001000100111101010000110101000000000000000101011101110001000000010011001100000101000001001111010101010100111101110100000100010100010101111101110000001111111101111111111101010001001101011101010001010001001101000101000011111100001100000100010000110100010000111100110011110100010011011100001100000111110100000100011100001100010011000000011100010101111100011101010101110000010000000111,512'b01000011111101000101000001110000010100010100010000010011111111000001000011110000010111001111010101010000010000000101000011010011110100001111001100110011110001111111011101000001000101111100110001010100010101110011000001000111001101010111110001001100010100010111110011000001010101110000010000000100010100010100110000111101001101000001111111011111010111110000011111010111110100001101111100000111110000001101000000001101001111111100001100010001000101110111110100010001010101110100000101011100111101000100010000110000,512'b01011101000100000001010000000011110011000101000101011111010101110000001100000111010000010101011101001101111111111100000000110101011100110100010000111101110001110011000100001111000000110011010101011100010011110001001101010000110011110011001100110111001101011101000011111100010011011100001100010001010101110011001111000101110111010000000111111100010100110001011101010000110111111100001101000101011100011100110001010101010100001101000100010111110000000100010001001111010100000101011111110100111111011101010000000011,512'b00010100010000111101111100001101111111010011000100110011110100000100111101110000110000000001011100000101110000001111010000110100110100010111010101000101110100111111110101000011000100110000000011000001110111001111000111000011000101111101011101010101000100010000001100010001011111001111010111010101110000001100001100111111001111011111011111000111000000000100010101110101011111010001110001001100011111111111110101010000000101110001000001000000011111110000011111010100000111011111000100011111001111110000010100000001,512'b01001100010100110001000101010111010000111111000100010101110000110011110000110100000111010001000101110011110011110000000011010101000001110111110001111111010001110000001101110001111100110111110101110000111111111100110011110000000000011111010111010011011100010000000000010011000101001100110000111101111101000011110000010011110011010100000111000011001111000101010000010100111111011101010000010001010001001100010001001101110100111111000001000111001100110000001111110101110001110001111100010100000111110111000101010001,512'b11110101010001110011000100001100010100110100110100001111010000001111000000010000010001000000111101010100010001000001000011001101110000010011010000110001110000010101011100010000001101011100001100011100001111110011110100001101010001011100110111000111010111110101001101000011111111000001000000001111011100111100000111010100001100010011110011111101000000010011111101010000001101010111111100001101000100000000000000110101000000010011110111111111010011110111111101111100110000111111001101111100011111001100000101000001,512'b00111100010011111101010001011100111111010001011111110101001111110100000100000000000111000000110111110111110011001100111111001111001100111101000001011111011100001101110011110111011111011101111101000101110000000000110001010001000011000000000111110001000011000011110000111111000011111111000011000111000101011111000100000100111101110111010001010111111101010000000101000000011100000101110000110001000101001100001101111111010100110111000100000100000111000001000001010001001100000101110000000001010101000100010001011100,512'b11011111010111011100000011001111011111000000001101111101010100000111011100010100010011000000110111010011000001111101110001110011011100010001000100110001010100011101000101010100011100110011111101110101010111001101001111000011001100010001000000111101110100010101111101011101111101010100110111010001110000111100001101001101110000110011011111110100110000110101011100010011010011010000000011000111111101000000010101000000000001110000111101010100111111001101111100110100010111011111001111011100011111000101010101010100,512'b00001100010101011101000011110101000101000100011101010011000100110000000000011101010001111100001100010100110000010000111111110001010001000011010011111101000101010111000101010101110100110100000111111111000001111100000001010100110111001111111101000000110100110100010100000000010100001100011101111111001111110100000001011101110000000000011100010001111100011100011101111101000000000000111101001101000100011111000001000000000000000101010000000111010000011100111100000000010001001111001111110101110100110100011101110000,512'b01110000010100110011011100010000010111011100011101000100110001110100000011000000010000000101010000010011000111011100000001001100010000010111000100001111111111010100011100111111010001000101000011011101110100000100010000110100010111001100010000111100000111110011110001010000010000110111010100000100000000000100110011110000000011110000000011000000001111001100010011110100000011001111000100000000110001010001110000001100000101110000011100110011110111110001010101000000001101001100110111010000010000110100110000010111,512'b11110000111111010000001100000000110111110011001111110000110001000011010111010100110101011101010001001100000011110011011111000011001100001100010001000001011111000100001111001101111100001100010011000011000001110101001100000100000000000100000011011100111101110100110011110000010001110100000001001101000000011111110001000111000100010101000000000001010111110001011111000001110100000001011101111111001111011100110101010101000100001111110101110011010111001111001100000100001100001101011100000111000111000100110100011101,512'b01110111011111010000111111010001000011000001001111010000110111010011000100011111000000110101010001111100000100000000001101010111110000001100001100111100001101111111000000010011000011111101000100111111010101110100111111110011000011001101000111000100011111000100001111110011111100111111000111111101111101010111001101010111110001110000000111001100011111110111010001000011000000010001110011010000000000110100110001010111010001110011001101000001001100011100110101011100111100011100111101110101110111010101110101001111,512'b11010100000001000101011101000011111100110100000000000001110001110000000101110100110011000001010011110000000001110111000100110000010101011111010001001100010000000000010001110000110100000100110101010000001100010011010011010000110001111101110000000100000100111101010100000011000001000111010000001100110111110011110011000001111111110101000000110011111111110000000111000000010011011101010101110000000100010001010000001101010101111101010100001101000101001100001101110000000101000100110001001100001111001100000100010001,512'b00110001000001010011010001110001000101000001001111001101010011110000010000110100001100110100001101110001001101110100010000010100000001110011010011001101111101000011000111000100111111000100111100000101001101011101010011000011001101001100011100111111011101000001000001110011010101000000000011000000010011110000111100000001111111010011011100000001110001010101000000001111000101001100000000110001001100001101110000110111001111010011011100011100001111111101111101011100011111011100111111111101011101110100110001110111,512'b01001100010011000000110100000011000100110001011100000101110101001101010111011100110000000011011100010001010101010100111111001100110100111100110111000111001101110001000111001101000011111100110000010111110011110100010000010001001101001100011111000000110000011100111101010100110100110000011111111100110000010001110000000100111111010000011101110111111100011111110100001101110011010011110000110000010001001101010011001100110001110000000100111101000001000111110111110001111111001101001100010000000000010001011101010001,512'b11011100010100011100000111110001010111111111110001000111000111000100010011010011011100111111001101000101010001110101010001110100000101110100000101010100000111000111110111011101000100001111001101000101110100000011000111111100000101010000000001000000000000000011110111010111000011010101000000001101111101010001110011000011011101010011010111010011110001000000011101010000000101001111011111010011001100000101110000000100111101011111011111000000001111010111010101000000000111000111010001010001000000011101010101001111,512'b00010101011101000011110111010111111111010011000001001100010000001100110001010001110111011111110000000000110011010011000011010111010001110100011101000100001101010111001100110000010100111100000011011100000100010011000100001111111100110000010000111101000101010111011101010100111100110100000101010001001111110001110111111100001100111101010000001111010001001101111101000011110111000100000001001101000111011100111111000100010001111111001111110101000001110101010111110100010101111100010000110000010011110011110001110001,512'b11110101010001110100011100001101110101001100000101000011110001111100011100110111110001000011000111010111000100010011010011001101010100000111010000110011110111010001111111011111010111110100110001111100000011010001111111011100110100000000110111000111011111011101110011010100010011111100010000000111010101110100110001000100010111000100010100011111110111110001110011111100110000010100011101111101000111111101000101110101111100110011111100110101110111000101000000000000010000000100000111001111011111000000000000000111,512'b01001100000011001101111111011111111101010100010111110000000011010011110000010001000100010011000101110111110011001101000000000101000100110011011101110001010101000100110011000111111100000001010001000001001100001111010011000100110011010111000100000000010001011100000100010101010011010011011101010100010000010111000001011101000111000101001111000001010001110011000000000101110100110000000001001111000111001100000101001101110000000000010101000011011101010011110111110101000000010001011100110000001111110000010100000000,512'b01110000000100000000010011011100110001000100010000001111010000110000000000010000001101010111110100001111010100010001000111010001001101010111010011111111010100110000000000110011001100110100010111000111001111000000110000001111000111110100011111110111010100110101001111011101001101000000010000011111010001011111110111110100000101111100010000110011111111001101010100001111000001000011000000000001000001110011000001001100000000110100010000111111110111000011000001001100010111110001000011110001001100111101110001110101,512'b11111100000011011101000011111101110001110111110100000000000100010000110011011111011101110001011111010000010111010001010000011100110101110100000111001100111100111101000011110101010111000011010000000111111100111100001100011101111100010000011101111100000001110011001101110000110011010000010011010000000111110100000111000000001100000111000111110100001100011100000101111101001101001111110100000011001101000000001100010000010111010101011100000001110101111101000011010011011100110100010111000011001111010000011111000011,512'b00110111111111001111011101110100111111110000110101110001111100000000110011111101000000001100001111000111011101000011001100011100110101010111000000001101000100000000110000111100010011110111000111001100001101110001111111110100111100110100110111000011000000011100010100001101000111111101010000010011110001000101010111010100110001000100001100010011000000111100110100000101010111011111000011111101111101111101011100000001010101001100111111010011000001000000011101010111110000010100000000010111010000000000011111000111,512'b01010000001101010000011111010111110000001100001101110011001101110000001100010011011100110001111101000000111100111100000100000100001111000001000001001100001101110000010011111111000101000111111101010000001100010011010100000001000011111111110111000011010000110111001101000001111100000000010111011100011101110100000011010000010101010000000000110001001111010111001100110001110000111111001111000011010011011111110111111101001111000111000000110011000100010000001111111100010100110011110111110000111101000111111101010011,512'b11010000000111010000000011111101010100000011000001110101110111011100110001110101000111110100000011000100000100110101111111110101111100000000000101001111011100010111110011000111110000000001110100110001011111110001000000110001010100010100001111000100011111000001001100110000001101110011111100000000011111111101110000000001000001110001010101001111000111010011110111110011010000000011000011001111110001110001110000000101010000000001110000110111110100010000110100011101011101011111110101000101001100010101011100111100,512'b00110011011100110011001101000001000011110111110111001101001111000011010111000100001101001101010100110101000011110011010011110001110000010011000101010011000111110000110111000111110001010111010011010000000111111101000011010011000011001100110011010000000100011111010001000000011111010111110101110011110011110101110000010111011101000001111111010011110000000100000111110101001111110100010000110100110000000011001100011111001111010000001101110101010101010011010100000000000100000011010000000111110011110111011100111100,512'b11110001110111111111011100111101001101000000111100011111110100110000011111010001011111001111010000110001110011010000110101011100000000000111000001010101010011010001000001000100001100010100010001000111011101110001110101011111010011110001011100110011010100011111111101111100111101110001000011111100001111111101000001111100110100011100000011010100011111000101010100110001010011000000011111010001110100000000011100110100010100010101010000000100000000000100011100001100010001010101110001111101111100010100111111000101,512'b11011111011111010011011100111111000111000011110000000001000100000011010001111100011101010001010011010100000101011100110011011101011100000011000111010111001100001101110100010100110001000000000111000111111101010100110011011101000000110011010101001101010011111111001111000001010011010111001100110000010000001100000001110001000101111100000100110011000000011101110011001101010001110111010000010001011100111100000011000101010011010100110111011100010100000001110001110001011101110111001100010000001101010011011100000000,512'b00111101000001110011010011001111010001011101010000011100011100011111010100000111000111111100010101000011000000111100110001000101000001001100001111010001001111010011110000010111110100010101110011111100110011110100010111001111000100011111000100010101000101001111010000010000000011110100010011000111110011010000000000011111110101110001000011110111010100000011000111001100000100010101001111110100000100011101011100010111010111110011011100000001111100000100000101000000110001000000010111010111110011001101110100000000,512'b01111101001101010011010000110001010000000001010111000001111101000101111111110111011111110001110111001100010011010100000001000111010101010000110100110100110000010001011101000011011100001111111100010000010100010101110001010101110011110100000100010001010100000001110001001111010100001100010101000011010000110100000000011100010111001101000100110101001100010101001111110000011111111100010101010000010100001111000001110111011111000001000011010011110111000111011111111100010001000100111100001101010100001111010100110101,512'b01110011010001000001001100000001010100111111001101010111111101111101010100000100000111000111010000010100011111110000110000001100010001110100000101010111111101111101110100111101110111000000110000011101000101000100111101000000011101010101000100110100000001000111110011011100110001110011010001111101001100000001000101000001010001010001001100110000110001000001111101110111011101111100010100001101010100001111010011000111111111011101010000010000010011000000011100110000110000010100110011110111000011111111110100010011,512'b00000100000011000000110011011100011101111101001101001111111101010111111100010111001111010101001111010111110000011100110111000101010001010000011100001100010111111100110101110100111100010000110001010011110111000101111100111111000001011100000000110111010101011111001111010100000011010001110100111101001100111100000011110100011100111101111100000000000011010000111101110000010101011111010100110101110000000101011111010100110101011101110011010101110000011111001111000000111100010000010001000101010011011111000011000101,512'b11111111000001000011011100010001110011111111111100000100010111011100001100000100001100110001110100011101001111111100001100000001001111010100010011110111001101000111000111001111010000000001110001000011011101011100111111110111110101010011010100010111001100110001000000110000010100111111110100001101110011111101110011010111000101111101000001110001110100010000001101110101010111110000001111110111010001110000111111001100010100111100010001010000110100111101000001110000000000000111010001110001000000010000010000000100,512'b01110111000001010101010001110000000100011101000011010100000111010100010111010000010101110001001100001100110000011100000001110001001111111100011111000111110001000000010101010100000100110111000000010000011101001111110011011100001100110000010001111101011111001111111111010011010000110000010011000111111101011111010111000101110100000001000011000011000000010011000100010100000001110111110100110001110000010000000000111111000111001111001111110000010011111100000101000011011100111100000011110101110001110001000000111100,512'b11001100110001010111000000000101110101010011000100000100110001010111110000000111110101001101000111000011000101000001000100111101000011011100011100011101010111110001111111110000110001110100010111000111000101110100000000010100000011010011001101010100110001111111110100001100110000111100111101110011010100111101000001110100001111010111001100011101000011110000000000000100010101111100110000000000110000111100010000001111010001010001001111001100000001001101011111001100000001111111110111000000010101110001110011000001,512'b00000111010000010101110111001101000100110100000101110111000100010111010000111100000100111100000000000111001100110101011111011111110011111101011100000011110001010101000001110111110111001100111100000000000100000111111111001101001100110001000000010000110001000111000011011111000000110111011111000001111100010101011100010111000100110000011100110100110011001100010001010100001100000101001111110100010000110111010000011111000001000000010000001111000000000000110000010100000011111101110001010111001101000000000011110000,512'b11011100110011001111110100110011000001000001010100010000000000110000110011110100010100000000111101010001111101001101010111011100110000110001110100000001110001111101000001011111011101110000000001000011111101010111010000110100111100010001110000001111000001110111110111001101111100000011010001011100011111010101010000000100000111110100000011010111010100001111010111010011010011111100111111001101110001110011110100110011011100011111001100111100001100110111010000001100000111110011110000010000011101000001001111000100,512'b00011101000001000100110100010111110100010101011111110101010100010011110000110111010011001100111100000101000000010001010111001101000101110100011111001111000000011111001111110011000100000100010000001100110101110000001100110001110111110100110011010111000111000111000011110000110001000111110101110011011101001100001101110011000011000100010001000101010001011100110101010111010011010101010100001100000011010011000011011101111101010000011101000111011101110111111111010101110000110111010111000101000000011101000001111100,512'b00011101000100110000111101110011010101111100000001010001011111111100001111000001000101000101001101000100110100110101000011000101110011010000110000001111111111001100111101110111001100000100000011110111001100010100111111000101110001011100010111111101000111000000000101000000000000000011110011001111001100000101011100110001010100000000110111110011000011110011001100110101110100010011011111110001000100001111000101110011000101110000110011000000011111110001111101001100001100000000000100110011000000011111010111011100,512'b11010001111100010001000111010000000100000101010000001101010111001101010100110001001101110001110101011100011100111100110011010001110011000001001111000011011100111111001101000001010001011100010100110111011100011101010111010011000001011100110100000101001100010101010011110001010011010001111111000011001100011111000011011111000011010000011101010101011101001101111101000111110100010111110001111101010100011100110000110001110000111101011101001111010000000000111100010111011100000001110011010111110000000000110101000001,512'b11110000010100000011000000010101000100010001111101001100010000010100010001001101110011001100110100001100001100110100010101000100111100110001110011011101000111010101000101010000011101010101011111110111000101000011010001010100110111010001011100010000010111010000111100000000000000000100111111110011000001010100001100110000011101010011010101010101111101011100000101110111000001111111000001000100010100011111110111000101001111111101011111000100000001110101011101010001010001010000111100011111000000000001000000010101,512'b00010000010011001101010001000011110000011111000001010011110100011111001100000000000001000100010111010001110111011101011100010100000000110011010101111111110000010011011111110100010100110000111101001101000111001101000101001101111111111100000000110101110101000001001111110100010011110011000101000111010111000000110000001111000101111101011101000000000011010001010011000001000001010011111111011100011111000001010001010100110101111100001101110100011100001111110011000000111101001101110000000100111100010000000011110001,512'b11001100010111001100011101000100110000011100000001111100001111011100000000111111001100000000010000000000000001010111011101110100010100001100000001001100111111011101111100011101001101000000001111011111011100011100000011110011000000011101001101000001010011110001010011011101110011110100010111010101000100000101000101000001111100000000010000110001111100001100110101000100010100010111110101010100001100001100010000011111110100110011000001010001110011111111111111110111000100010000110100010001000101000011011100110000,512'b01001100010111010111010111010001000000001101000111110000010000000011011101011101110011000111000011000011010100010100000000010000011100001100010001000100110011000101000100110000000100001100010100001100000000111100110011000001000101000001000000000001000000010101000000000101111101110011110111110011110001110011010001010011111111111111001100001100010001010001000001011100000001010100110101111100010001001111000001000100110101110001000001110111010011010100010101001101000000000011000100011111010011000001010111111100,512'b11110001000011010011110000000101000100000111110000110100000000010100000000001111011100000001111100010011000000001111000000010001110001111111000101110000110011000000010011010111001101010001000100111111010011001100010000000100110001111101000001110001001100110111001100010111111111001101000100111101010011011100000001000001010011010101000000010100111111110111010000110011010111000101000011001101010101110011000100110001111111000101110101000101000100010100111101000011000101000100110011011100011100011100110001010011,512'b01001101010111000100000101110011110000000011001101000011001100110001000100111101010111010000000001110101010000000001001101011101011111011100010101110001011111011100011100011101000001000001010111001101010000000011000101110001111100110111110000110100010101010111001100110011010001010000110000111111111101111111110000000100011101011100010100000011011111011101110011010011010001000000110101010101011101000111110100001101110100110100011101000001001100110001000101010001110101110001111111011100110100110100111100010001,512'b00000011010001000111001100000111110111010100001101010101010011001100111111011101001111110111010000010111111101001100000011110100000001000111000101110000111101000000010100010100000101110011110111110111110000111100010000111100010101010001000001110100110111010001011101010011000101000011000011010011010001110001000011011101111100001100111100011111110100001101110000010011001111110011000111010101010001111101011111011111000011001111011111010100011100010001011111001111110011010011001111111111000100001101011111011111,512'b00110000010000000001010100010000010011010111000001010011000100110001000111001111010100110111000011000100111101010011000101010000110000000011000011010111001111111101110100000100110000011101000000010101110000001101110101000100110100000101110001110001000011111101111101110111001111000000110000000101110101001111110100111100001100001100001101000011000001010001010000010011010101110011000101000111111101000000010011001101011101001101110001001100010011110100000001001111001111001100001111011111000101011100000100110101,512'b01010101000000011100010001011101010100001100010000110001000111110111001101010100000000111100010101000101000011010000111100010011000000000001110001000011000000010111110000000001011100011100010011110000010001000100110101000011000000010000000011010011110101011111011100110011010001001101000000000100011100010101110011000100001111000100001100010000110011011100010100110100110011011111000100000000000000000100010101000001010000010100010100000001111111010101011111000100110011001101010100000001000111000100010001111111,512'b00011111110101111101011111110101000001000100111100010111001100010100000100110011000011110001111101010011111100111101000100000100000100000100010111000000000001110100111100000111001100000001000011001101000001000100001101010001011100001111111101110101010001110000000001000000111101110011000000010000011111010000111101001101000001010100011101010100010001010000010101000101010100010011000011000011010000110011011101110111010001000000111100001101000111110111010100000100110011010011010101010011001111011100011111000100,512'b00110000000001110000111101001111110101001101000100000100111111001111110111111101000100111101000011010100011111010011000100000111010100010000000000010100110011011101111101010011010000000011000001110011110101010111111101011101111111011111010011000001011101110111010111010011011100110011010011000100000111011111010100000000001101111101000000001101010111000001001100110100010011000000110101000101110011001111010100000011010111001101000111110101000100000011001100110111000000000001111111001111001101110111111100001111,512'b11110011110101000100000000110111011111110111010100000011010111000100000001110101110111000000110111000011000100001111111101000011000100010000110001001101000001001101001101000011010011010111010111111101001100010000001100000001000111001101110011000000110011110000000001110001000011000111000011000111111100001101010111110001011111000101111100010111010001000011000111010101001100001100000011010001010001010101000000011101000101110111011100001100110000000111011111001100001101111111011111010101010011000011111111111101,512'b11010000111100010100000011000001111111111100011111110011001111010001010111010001010100000111000100000000110011001100000100010011110111000000110011010000000000111111110011110011110011010100001100111111110000111100010100010111010001010111010011110111001100000011010001000111000000110001001111000011000111000111001111011100000100110000010101001101000011011100011111111101000111000101000100011100001101000001110100010001011101011101000001000011111100011111110001001101010000010001010100011100000011001101010011010001,512'b00010001110011010111010000010000000000000011000111111111000000110101000100110001010111111111000000110001110001111100000111111101110100000000011101010101111111010111000000011111000000110100111101110000000011011100110011010001000000010011011101110111110111011101010011010000001100110111010111010000011101111100110001110111000000111111001111111100110001110000010101110100001111110111000011000000110000110111001111010011010100011111110000011111110001010100000011010101110001000011000001000000010011110000110000000001,512'b01010100010111000100111100011100000000110100010001010101000000110101011100111101110101111100010001010111111100010111001100110111001100110000000011000111110000000100111111010111000100000011010000110001011111001100010101010000000101010000000000010101010000000000000111001101000011000100000101110011010011010111001100110101001101010001110000010011110011000000011100001100010011010000110001111100000100000000000001110011010001111101010111000000010100010011110001110101001100010011011101111111011100000000110000010001,512'b01010001000011010001110000000000000011110111000001011100011111010011110111001100001100010011000000110100110011000000000000000000000100110100010001010000000011010101110001111100110011010011011101110011010100110001000100001101110100010001110100010011010000011111010011010111011101010000000001110001010011010000011111000000110101000011000011111111001100001111010100000000000101110101111100001100001111010011110000110001010011010001001111111100000001001100110100111100110111010000011101001111010111000101000101110100,512'b00010100110011110111110111111101001101110000000001010101001101001111110011111111010001010111000000000101011101001111001100111101000111000111110100011111110000110101011101011101111101110011001111000100111101110000110001000000110000010111111100000001000001010100000000010101010100111111000000001100000011110101110100011111110001000100010001001100110101000100111101000000011100111100010100111101000000000100111100000001111111011111111111000011110100000111000000110001000001010101110000111101000001010000001111111101,512'b11011100000111000000000001000011110011000100001100110001010000010011010101010100010001000001110111000111000101001100010111001111010000000101111100110100000001010100000011011111001101011101010111011111000111110100111111111100001111010000011101010000000000010000110111001100000100000111000000010001000100110000010011110000010100000000010011110100110011010011000111000100010111011101000100010011110111010100110111010000000000000101000100111100011111010000111101111101110001011101111100110000000101110000111111010111,512'b01111101001100010100010000110111000101010101110100001111010001000100001111110101001100010000010011000000010101111101010011111100110101011100110011110011001111011101000001111111111101010101011111010000111100000011001111010001110111001111001111011100001101010100111100110100000011000000011100001100000100000011011100000011110100000100000001000001001101000001000000110000000111000001011100011101110000110000010000010111010011110111000011110000010001000000000111110100111100000001110001010001000100110000000100010011,512'b01110001000001000001011101010000000011000101111100110100000001010111010000110100111101111100010100110000010011010111000011000111110000110001111101011111000011010101110111110000110011001101111101000101110000010001000000001101000100010100011111010101110001001111110011110000110000001111010011000111110001110111010000011111011100011111010100000011010000001101001111000011000000110001001111011111011111010001010011110000110001111100000111010011001100010100000100011100000001000101000111000101010000000001110011010001,512'b11000000011111011100110100010011010101010101110101110111110011010111110000001101010111110000111111000101010000000001110000111100010001000100000000011100001101110001010101010001000101000000110001111101110001010011111101010001000101000011000000000100000111110001000101110000001100110111000101001100010101010001010100010101001100010100011100110111011101001111000100000001010011000001111101111111001100010000110111001100011111010000000000000111111111000001110101000011011101011101011101001100010101000011011101110011,512'b01000000110000011101000000110100110100010000010000000111000011010101111111001100010111000001010000010111011100111100110001011101110100010011110000000101000000010011011111110011000101110001010000110111110000001101000011010101000011011100000001001101011100110111000000011111110000010111001100110000000100110100001111111101001111110100010000010011110000110100001101110000001100010111000001000100110100110000000100110111011100000001110001000011001111010001000100010111111111110111110111110101010100000100010111001100,512'b00000011111111010100010111110000110011110011001100001100001111000000110011010001000011001101000001000000001111110100010101110011010101000001010011110111110111000001001101000100111111010011001100000011000011000100011101110001111100000000001100111101110001010001000001011101000000010111110101011111110000011111010100110101000001111101001100000000110100001100000101010100000011011101011111111111000000010011010000110000011101010000010011000101000000110000110100111100001100011111110000010100111111111100001101001111,512'b11110011010100110011000111111100110011001100010000110001110100000011010011001101010111000000110000010001110111000011010001111111000000111111000101111100011101010000001100000000111111010001110100011101110000110000000000000111000101011111000011110000010001110000111111001101010011110011110000110000110001000100110001010101000000110100000100010100001101000011000111011100000001010001000001110000110111000100011100010101110011110001110000110011000001010111110001000000010011011101011101011101000000000111010000110111,512'b01110011000011010101000000000101111100001101001111110101111111000001001100010001010100111111001100011101110000000000010111000100010011010001011101000001010100011111000001010011011101110101011100010001010000010101111111000101010000011100000011110111011101110000000100010001110011110011000001111100010011000011110000000000001101011111011101000000000111010001000100111101000000000100001111000100110111000100010000000001010000110001011111000100010100110100000101110011011101010000110011001100110000110100111100000100,512'b00110100010000000011010001010101000001000000000000010100110011001101111100110011011101011111010100011101110100011111010011010011011100010000001101000001000100010001000000000000000011001101110100111111001111011111000000001101010111010011000101010101010101010000000011000001001100000001010001011100010011111101001100110011010001010100010011011100111100110101010011111111111101010011110000011100111111000100110000000100010001000011001111011100000000010101110001110101001100010100011100000001111100000011010011111111,512'b11000101000101001111000101111111111100011101110100010100011101111101010000001100110011000000010000010001000100000100010000010011010000111101111100010011110101000011111100110000000011001101011100110100010000011100000101111101000000010101111111111101110011010111010000000000011100110100010001010000010000111111110011011101000000000001110001000100110000000000010000001111110101001100011100111111010100001101000011001101110011000000000111110000111111011100001100000011000101110111111111000000110111010001010111010101,512'b01110111010001000011000001011100000011001111110011010001010100000000010011000000111111011100000111010111000100000111000001001111010000010111111100010000010101010100001101001100111100110111110111000000111100000111000100110100111100010000000001000011000000111111011100010011010100110111110101110000000100010000000000000101111111000101110101000001000111110011001100110111001100111101000111001100010100110100110000111101000000110100111100111100011100010001110100000001010001000001001100010011010011000001000101111101,512'b00111101000001001101011100010011000101110001011101111111001111000000010101011101010001110100010000001111000101010001010100011111010011110101001101010001110100010000110111001101010100001111000001010000000100000111010100000101001111000011000100010100000101011100001100110011110001000100001111010100010011010000010111000101110001110000001101001111110011110011000011001111000001010011110011010011000001000000001100010101111100110111110000010011110001001101000000110100111101110011000011000011010001000001000101000100,512'b01001111110011000101110011010001001100000101011100110000010111011101000000000000000001000111000111010001110000000100110011001100011100011100110001010001110001001101001111000000011101110100110000010111110000010100010100010111010011011100010100010001110101011100010000010100000100111101110011000100010011110100110001001101110100000011011111010011111101000101000011110111000001110011010000000111011101000100001111011100010001010011010100110101000001000011111100000101010100110111011101011111110011011111110000110101,512'b11011111010011110011000011111100000000010001111111110011110011000101010000110011110101000000010101110000000011010000110101111101010001000101111101110011011111001101000111010100110000010001001100110100111101110111111101011111110101110011000111110000010101011101110000010100110000000000000000011101000000011101010000010001000100001101110000000101110011111100001111000000011111110011011111000000001111010111110111011111000101011101010111110000001100110101010000011111001100110111010011110000000011000001000101110001,512'b01000011001101111100000001111100010001110111011100011111000001000001000100111111001101110011001100001111111100000101000100000001000000110111110001010101110000010000110001110001001101011100111100111100110101001111010100000011011101010001010001011101011101000101001101010101001101010101000100110000011100000111010101111101110111000001110101111101000111001101110100110011001111111111111111000011001111011100000000000011010111001100000001010001010101110100000101000111111101000011001101011111010101111100110111011111,512'b01110000011100110011110000011111001111010101010101110011000001001101011101010100001100011100011111010001110000001101000011001111010001111100110111000100000011010100110001000001111111000100000111000001000011000111000011111101010000111101111101110111111111110101110111000001111100011100010000000111110001010011000000110101110101010001110011001101110000011111111100000011110001110011001111110011110111010000000000011100110000110001000111111100010011111111011100010111010111111100000111000101110000011100110111110100,512'b11001101110000010000001111001100010001001111000111010000110011110100010101001111110001010001000101000111110011000100010111000011000100001111000000010001110000000111000111010001000100000000000000010011111101111111110001000101000100010011110001010000010111010001000111010011110011110001010011011100110101000001010100000000001100111111011111110100000011011101110011110101110101010011110000010001011101001111001100000100001101010001000101000100010001001111110000000000001100010011010001110001010011011101110101010000,512'b11110111110111000100110000000011011111001111111111010001010011000011000100000101110000111111001100011111001100011101001100110000001100001100000011110011111101011101000011000000001111111100000101010001011101001101010011001100010001011100110100110101111101010000110000000000110100000011110101111101010000011111111111111101000001011111111101000000010100011100110001110111001100110001011100110101110001111101000011000000010011110101010111110011110011011101000101000000111101110111000100010001000101000101011100110101,512'b00010011000101110000110000000011110000111100111101111101010101111111000000010011000000000111000011011101110100010011010011110101111111010000110000010001010000010001011111110001000000111111110000001111010011010111110011010101010011001101011100110100111101110011001111001101110000110011000100011111011100010000010111010011110011110001000011011101010111110001001101010100000101110011000011010101111111011100110001110100000000110001110011111100001101010000010011011101001100010100011100111100000101010100010001000101,512'b11010000111100011101010111000000000000001100000101001111001111001111001111010000000000001111000111010000000000001101110000110101000000000111000000111100000111110100111111011101010001000100111111111111010001110000110011110011110001001100010111010101010001110011110001111111110001000100110100000000010101110100110100110101001111110011010000010101111100010101000011001111000000011101110111010111010011110001000101111111010100001111000101010000000000110111011101001101010001110100010011000101000000111100000001010011,512'b00000000111111110100000011110100010011001100001101000100010101011101010000110000011111010101000101110111111101011100010001001100111111010000010000010000010001110001110001001111000111010101001111000111010001000101000011011111010000001101010011010000110011110101110001000101010001001101010111110011000001010000110101000111010111000001010001000001000111110101011100110000011101110100010100010011000001010011000001111111001100111111000101000111110100010011010000000011001100000100011100000011110000111100000000010100,512'b11010011010001110100011111000100010000110000000011001100110000010100110001001100001101011111000101011101000100110011010011110111000111111101110000001111000001000011110101000100111111010011011100110001110100011100010000000001000000010100111111110000110101010100010001011111111111010111110001111111000100110000110000110011000001001100110101001101010100000100110100000100000101000001111100011100110100000000110111011111000111000111000011000011011100110101001111011111001100000100010000000111000100111101011100011100,512'b01110001001101010011111101010000010101110000010111000111000001110000110111010000010000010000011100011100000100010100110000111111110100110100000100010111000001000011011101110000000000010100010000010101000011000000110101001111000000010111000001000000110100000000000001001101011100011100000111000001110111000000010101111111001100000001010011001100110101011101010000001100011101000100011111010100000100001100110001010000110100110001111101001101110111010111011100010111000111111101110011011111110001010011010011000111,512'b00000111000100000000001100001111110011011111000011001101000000110011000001110001000000000001000101011101001100000101010011011111001101010001000011000100000000110101010100010101110011111101001111010111010100001111110000000000010000010100110101110101000101011101110000010011110111000100000001010100110100001100000100110100001100000011000100110000110011111100000100001111000101000101000111110000000000010001110111010011000001010000010000001111000111000001000001011101000111111111110000111101111100000001110011111100,512'b01010111000100000000111100010001000101001111000100000011000100110111000011110111001100010100010011000001110001001100010111110011000001000001001111111101111101010000001101010100001111000100010001000000011111110111110111110100010011000000000100110011110101010000110100000001111101000000110011000000111100010011010101000011000011001100000101010001001101110000110111111111011101010100111101000011110001000111111111010111110100110111000001010100010100110011010101111100011100001100000001011101000000110011011101010100,512'b01011101010101110000110111000111010101011111011111010111010100010100010100010111110000010101110000010000110011001101010000110111010011110000110111110100110000111101000101001111001100110111001111111100001111111101000011010011110100000100000100011101001111010000011101110000010011001100111101001101000000110111010011000101011100010001001101010100000101000000111111010001001111000111001111010111010001001101110011000011110000000011011101000000001111011111000101000011000001000001110000001101000011000100000001011100,512'b00110011000000010101010001010011010001110000000001001100010101000101010000000011111100001100010101001111111111010101000001010000000000010111010000010001011101110100000001110111010001110001010000000101010101110001110001010011011100000000010000011100010100111111000100010001000011000111010101111100011111010001000000010100000111011100010001110101001101000011110000110111011111001111011111010001010011110111110000010000000101111101001111000111010000111111110000000111000000010100110001000000010001111101011101000100,512'b00011101010011010000010011111100010100110111111100000101010001010011000000110101000011111101010111000101111100001100111100001111001100111100110111111111001111010100110011111100110000000101011111111111110000000100001101001111000000011101010111010011110000010100000101110101000100111101000100011100110111110000000111001111110101010011000011110011010101001101000011111111000100000011010011000100000000011111001101111100001100110000000101000000000000010111110001000100010011010100000001010101110101110000110100000100,512'b00010101010100000101010111110111000101010111111100010011010111000000011100010100110000111101010100111100110000010011000111110100010001001100110011000000110101010111011100110001111101001111010100111111010000110001000011000011011101110101010001001101001100000000000001010100000000010111110100111100010000000111010000110011000111000001011100110000111100111100011100011100011111010011000101001101011101010100000101110111111111110111001100000100000101110100010011110000000000000100001101001100000101000000000111011100,512'b01110100000000110001110000110000010101110100000000111111000011011111110000111111001101010011111100000111000100111101001111110001110000000111111111000000010100111111000100110111000111000000001101010011000100000001110000010011110000110011001100000101111101000111000000010011010000000100000100111111000001011101000000111111111101010000111100000001010100010100010101110101000100010100111111000001000011110011111111001101110000011111111100000000110011110001111111110111110011010100010100011111000000111111001101011100,512'b11001100010011010001000111110000001111110001110001010111000100000111010000010000110001010000010000110001110011001111010001001111010101000011010100001101111100011111110000010001010111001100010001011100010001110100111111110011010001001111001111001111010111001101110101111100000011001100111100110111010111110101010011110000110100111111110000001111111111000111010111000111110111001111111100110111110111010000000111110011000100000011001111110100000101011111110111000100110001011101000001110101110000110101000000011111,512'b01001111001111010000000100010000000100110000000011111100110100110011001111011101001101000101110001011101000100011100111101001101111100001100110000000011010111000111011111000101001100000100000011110001010101000100001100010001010001000001010001001100110011110100001111000111110101000100000101010111111111000000000111011111000000110100110001010100001100110011001100010101001100000001001111111101001111001111110011000000001101010101010001000001110100111100010011001111000101111100010001011111001100010011000100000100,512'b00110011000111000011010001010011111111010011001111000011110111011100111100011101010000000101010011110000110001000100010100000011000100110101111100110011110011000000000000000001110101010100001101111100000000001100000011010001010001011111010101001111110001000100010001010100000111000011001111000100110100111111000101000111111101011100000100110101010001000001110000001111001101110111010111001100000000000001010101010100110011010000110000111101111100001111111100111111010001010000110011110001110111010000111101110001,512'b01000111110101001100000100110011111111000000000111001100011101110000110111110011011101000111110001001111011100010011111100000111010000011100110101010111000000110100110000011100000001000001110100000011000100001100111101000100000100010000001101110100110011010101011111000101010000110100000100110011111100010011011101001100000000110011000100010101001100110000111100110001011101110100111100010000010100000000000001000101110101010000010000000001111100011100010111001101010011110100000000010011000000110011110000000101,512'b11000000000101111101001100010100011111110011011100001101000111010000010000111100011100000111110000110011001100000011110100010000001100001100010100000011110000110000110001110100010001010100001100000111110011000100010001000111001111000111010100010001110100011100001101110111010000110001010101111100001100001111110000001100001111010011110100011100000000000000111100111100000000000101011101010011000000000011000011000101011100010111011111110011110001000111111101110001011100011111011101010001001101000111110000000101,512'b01000111110000001101011101000000011100000011110000000100010101000101010111010101111100010011001101011100110100010000000101010001000100001101010111010001001100110000111100110001110001110000001101001101110011110101010001001100010100110001111111001101000000110000110111000101001111010101010100010011000001010000111101110100000111010001000001000100110101000011000000001101110111011101110000000100010111111100010000110000111101111100000111001100001100010011001111001101001100000001110101110111110001000000011111011100,512'b11010001001100000101010001000011110100011101011100000001010001001101111100110100000000000111110011011111000101110001110000000100110111001100110100110011000000111111110001110001010101000101001111110111000011010100010100110001110000000100010001001100011111000000111100011111110100000100000101010100000011000001010101000011110001001101011111000101001100000011000000000000110000000000001101000000111101000100111111110000111111010101001100010000001111011101110001011100000000001101010100110101010000110100110101010101,512'b01000001000111111100000101000011010011110011010101000001010100110000010000010100110000010011000001110100000001110000001100110001000100110000001111010011011111000011111101010100000001010011001111000011001111000001010001001100110000110100111111001111000001111100001100000000000001111111000001010100010000001101011100000111110101000001000100110111000111110100111111110001001101001100011111010101010011110001000001010000000101010011011111111111000100110100111101010000000001000101110001011100011111000100011111001100,512'b00000101001100110000110000000111001100011101000101001111011100110011000101011101110101111101110000010100000101111111000011110000011100010001010000000111011100000100000011111100010000000011011100110001110000010011000000010111001111110100110101000001110000011101110000010101110000000000001111110111110000111111000001000000001100000001000000010001010001001101111100111101110111010011000011111100110000000001110011010101000101110001010001011101010001000111111111010101001111011111000011010001010000010101001100011100,512'b00001100000111110011110001111111000000000011011101110000000011111101000000110101010101000111111100000100010011000000000100000001110000001101010001010101000100000011010011001101001100010001001101000100000100110011011111000111000100011100011101010001000011000001010100000111010011000101010011011100010100110011011100000100000000001100011111110000001101011101000111010000001111010100110100110011011100110101110011001111011101010101111100110001000000010100110100000000000100000001110001011111111101011100011111110000,512'b11010000001111010001000000000001010000010000000001010100001111111101000101010000010001010011110000010111011111110100110100110101010100010111001101001101000111010001110011010111010000000000001101111100110001001101001101110001110100011100010101010000000111000001010000000101010100111100010001110111110000010011110101001100000101011100110100111100011100011101110111110101110000011101000000010100001111001101000011000100000000010011110011110001110101111101000001110011001111000101000000010100000001111101001101000101,512'b11010001110111000100000011000011001101110001001111011111000001111111000011011100111100010011010101010000000100110101001101110100110000000111001101001100001100110000110101000111010100110000111100000000010000111101010011111100110001010011000101011111000000010011111101110111010000110111000011000011110100000000010000010100010111110111010000010111110100111100010011000111011111000101110011111100001101000001110000011100111101000001110100010011000100000000111111010111110001110101110011110000010011000100000100011101,512'b11001101010011110100111100111101000111111100010101010000110111111111011101111111010011001101110101111111000001110011000011110000111101010011000101001100000100001111000100110011111111000001000001011111010001000101001101110011010100010101010011010011000101110100000001110011110100010000110000011101000001010000001100000101011111001101001101010011010011010001010111011101001100001101001111010101010001001111110001000001110100001101011100111101011100010101001111011111001100000111110100110111010001001100010111110001,512'b00011100110001111101111100110100111101001100110001001101111101010011110000110000010001001101010111000011011100000000011101110111011111000101010001000000000011000011010111011100001101111100011100110011111111001101000111110001111111000101000100011100010100000000110100010000011111110011111111110001001111000000010001000001010000000101110011001111000000110101000100000001111111000101011100111100010001000001110111000000010001010001001100110011010111000101001100000101010111000101000100000011111100010000010100111111,512'b00110101010000010100111111111100010000011111110011010000110111010001001111110001110011110111110000000111010011010001000101000101010000001100001101000001110011000101011100000011000001011101010101110101111111000000110100000111000100110100111100010101000001011111001100110001110011000101001101010000001101001100011100110111000111000100111100111100001101011111001100110101010000110111000000110001111101001111111100010011011111010000110011110111111100110111111100110111010101011111000011110101110111010000010100010000,512'b11011101001100000111110001010111010001011101010101011111000000110001010000000000110100010001000001110000110111110000000000000111000111110101110000000011000011000111000001000001000100001111110111000101000011000111110101000111000001000111010111000101010000000111010011110000000001011111011101001101001111000000011111001100000111010101011101000100000011010000110101010001011101010111000111110001000100001111110011000100000001001111110100110011110101110001111101110011111111110001010100010111000011111100000100001111,512'b11000000000111111100001100000100010100000000010000010000110100110001000000111100011111010000010000000000110100110111110101110101111100111100001111010000110001000100110001000101000000010011010111110001000000110011110011010111010101011100111100110000010111110001111100000000010100111101111101110000000000010011010000010111110100011111110101010011010000111111000101010100010011111100010111000001010011110100000011110001000011011111001100011100110001001111010000111100000000000001110001110100000100011111010111000111,512'b00001101110001010001010011110001011100000111000000000111110001001100110011110101011100110101000000110101000100110001010101110111110111010000000101110101010001001101000011010100111100010000110100010000011111010001110000111100110111110011010001000100010100000001001111000001010100000111010011011101000101110011110000011100111111000100110011000100110000010001110011111100110100001111001100011100110100000000000000110001110101000101110001110011110100110011000101000001010111001111001100110101011111011100110000000011,512'b01000011011101011101111100000000110111011111000101110101110011011101011100110100000011110001000000001111010111010111001100110011010101110101010011010100111100000011011101111111000100111100010000111100110111111100110101001101000101010001000011110111011111000000110101000100011111000000000001000111000111110101000101001100010100000011001111111100000111000101110100001111000100010111110001110000000111110011000000010000010100000111000000011111000100110100010011010000000000000100011101000011011100110001111100010101,512'b00111111000001001111000111010000010111010000111100110101000000111100000100001101110000110111110000011100010100001111011101110101010100001100110001010101010111110111010100011101110001001101000011111101110001110101000011111100011111000111010011111100010011111101110101110101010111010100011100000011001100011111110111000011011111010001111101001111010011010100111100110000110100011111011100110111011100011101011101111111001100010101111111110001010100010001000000001111010011000001110000000000010100010001111111110011,512'b00000000001100001100000001000100110111111111110100010111111111010001000011001111011101000011010001000101111111000000010011011111010000010000110000001100111100111100010000110000000100010000111100110001011100011111001111000100000100000011110101110100110000001100011100110100111100010000011111111100110000001100000011010101010001110111010001001100010101001111111100110100010101000000010001000011111111110000000000010100010001111111001111011100000101011101110100000111110111110000001100000101111100010101011101010001,512'b00000100000101010100010000011111000001111111010100110101011101111101110001001100110101111101010000010111010000111100000011110011110011010011010111111111000011000101000101111101000111110101010101000000000111001100010011011111000100010111110011011100010100111111010000010100011100010001111101000011000000010001001100110011111111110000011111110001011100000001111101000011001111001111000000110001111100000100010100000000010001111100010000110001111111011101001100001100110001010000111101001101001111000111000001110011,512'b01011101010101000011010000000101001111000101000011010101001100110100110001000011000100001111110100111101000000000111111111011101110000010000001100000111110000111111111111000100010101000100010001010001001101000001110011000100001100001101001111011101110111011100001100000001000011000101000001110001111100110100010011111100000001000100000101010101110101110000010100010011110000001100000011111111010111001100000101110000111100010000001100111101010001001101110111010100000000110000011101010111010100000001110000010001,512'b11110111111100111111010100000100000100111111111100110100000101010100001111110100110101001111010101001101110111011100110011010001000100110001110000010001000001110101000100000011000100010011000001000111110100011111111100011100010111011100110111001101110011110111000000010001000111001111011101000001010011111101000111000100001111010001001101000000110111010011010001010111000011111111011101110101001101110011000101010111110000000111010011000001001100110000001101110000010111110011111100000011110111000001000011110100,512'b00000000000000110111010101010000011101010011011111000111011111001101000000001111010000000001110000010111110101000100110101110000000001110001000001111111010000010100001101011111000100110111001101010011000111010001011100011101010111000001110111000001001100000000010000111111010100011100010011010000000000110100000001000101000111110000001100000100010000000000111101001101110101000100011100110100010011000011110100000111001101000000111111000001010111000101110000010000000001110111001111111100011100010011011111011100,512'b00110100011100111111110000000000111101001101000011000111000001010000010011000001000001001100000101000100110000111101010111010111111101111101110011011111010011000100010001000100110100010100000111001111110111000000110001000001110000010011110100001100011111000000011111001100110111000011001101110011000000111100110001000111111101000011001101010111110101000001010011110011010101110111000011110100010001110111001100010100000101011100000100000101010000000111111100110000111100011100000101010111000111010011000000000000,512'b01010100000100001111001101110101000001111100000111010100110001011101111101001111011101011101011111110111111111110000010101111101000001110111000000010011010111000111110011000111110001000001000111011100011100000011110100111100001101000100001111011100000101110101111100010011010100001100110011000001000000011100001101001100011111000111011101010100000011010111000111000100000100111101001101000001110000000111001100011100001100000001010000111111001100110001011101000000001101000101010100110111110011111111111100110100,512'b00111100000100000100110111000011110001000111000011010100110111110100110011111100000101010101000000110000000100011100110001010001110000001111110011110111010100000011000001010000010000011111110011010111001111010100110101010111111111000111001101000101010011000001010000111111011100010000110001111100001101110111110100011100010001010011000100010001010111111101000100000100010111000101000100000001110000110001001111110100000101000000000011000011000011001100000101001100010001000101011100110001000000001111110100000000,512'b00110011111100000001011111000111110000001101000101111111010101000011001100010000001100010000110000111101010111001101110011110011001111111100000111111101001100010001000100001100111101010111010011110000010100111111000011110011001111000111111111010011011111000001000011000011110111010101110101010001111100010000010101110011111100111100110011010111010001110111000011000011010000000101000001011101000000001100110001011100010011000011000011010000000000000111010111000011010000110000001111110111010001001100011100111111,512'b11000000110001001111001111110111000100110011110111010101001111000100110011010000111100001101000101010000000111010011000101111111110011111101110111011111111101001100000000000011010000000011000000001111001101000111000111000100010101111111110100110111110011010011000100000011010100001101010001011100001100110000000101000101110001111100010100000100011111011100110100110111000011111100010111000101000001011100011100010011010000010000011100011111001100010011110101110001001100010011001100000111010111001100000100000100,512'b11010111000000000100010111010111001100001111111111000000110100111100010001110011011111011100111101011101001100000001110100001111000111010000001101110000000111010011000100001100111111010001000011001111000011000101000100110011010101110111001101011101000000000111010100000011010111110101110100001100001101001111011111010100001101111100011100110100011101110011000101111100010111000011111100011111011100001111000011000011011111111100001111110001111100010100011111000101000100001100010001011100010011110100110000001101,512'b01011101010001000000000001011101010111000000001101011100001111011101011100110100110101000101010111000100110111011101110000001100000101110011000011000100010100011111010001001101001111111100011101000111010011110111111101010000011101110001010101010000010000110011000011011100000101110101110001111111010011000011110001001100010011111100010000010001110001110100000011000100001100010011011111000100110011110101110001001100110101110001110000010011110111000001000100111100011111110011111111010011110000011100010011011111,512'b01000101010101010101110100000100011100010101000000010101011100010101110011110011010011110111010100110001001101110100110100011100110100000000010100011100000000010000110000000000001101011101000001000111010000000011010100000100110000011111110011001101010101000000010101000111010000010000110100110000111100110100000111010000110111000011110000110111000100111111110111110000010100001111111100000100010100110000110101011100110011110011000000010111010001001111110111011111011111011111000111000011110111001100110111010100,512'b01111101110100111101000000110011010101001100111100010000110111000100110001110111010100011111010111000011001101110111010111001111110111011101010001001100000000111100000111011100011111110100111100010011001111111100110100000001011111000101110100011111001111011111110011000000001101110100000011000101010011000101110100110011010011110111000100001100110000000111111111110101110011110111000011000011000011011100010000000000110001000100110101110101010111000101000000111101000000011111010111110101010000001111111111110011,512'b11010101000011000100001101010011110111010001000100010011010001010011011111110100010011000101111111110000010000000101000011010111000001111111011111010011000111001111011111001111010011010111110011000001011100000000110001110100011111011111110001010000110001110101110000110001000100011100110000110011000001010000110101110100001111000011110100010111001111010001010111000100001100110100000011000100111100001100010011000111111100000000110001011111010000000100000011011101110111000111000101110001001100001100110000110111,512'b00110000001100000111010000010011001111001101010111000011011111110111001100010001010001110001110001001100000000010100000000000111001101000100111100010000000111011100000000000111111100010100000000010011011111000111110000110001000011010111000111000100010100110001000111010000001101001101010000001111010100001100010000111101111100001111010100001101110111111111111100001100000000000000010100010100000000011101000111111100001100001100010001000011000100111111001111010101011100110100001100000000010000110000001100010100,512'b11000111111101110100000111000000110100111101010000011100011100111111000000110001010101010011000000010101111100010111111100111111110011001100000011000000110100011100000001000100000100110011000100111101001111000001000001000011000001110000010100000101011111000111010001010100000101011101110000000001110100011100110000000100110001111111110001111111111111010101010011010000110111110101000101111100000000000001001101000011000100000111011101000100001100110011011101111101110011000000000000001101000001110100000011010111,512'b01111100111101010000000111000000110000001101011111010100011100000001110101000100110001000011111101010101010100110101110000000011011100000100010100111101001111001100000100000111110100000111000101011111110000010100001111010101010111110000001101110011010101000000110101111100001111000100110011010000000011000000110101110101010100010011011101001100001111110111000111110000111101110001000111010001000100110011000101010011000011110001010111010011011101110101011100011111010011111111000000010001011101010000000111000111,512'b00000101010011000111110100111101010001110111000000111100001101000000010001011101001101000111110001110111000101110100000100110001010111010101000101110001001100011100010011000101110100000101010100001101000000011101110101110001110100010001000111000001111100110001000111111101000100000000000111001111001100110101000011110001110111010011010100001101001101011101010101010011000100001111001100110001010100000001010011110111010101111111000001001111010100001111000001110111010101111111111100000001000000110111011111000000,512'b00010011111101111100010000110100011100000001001101110100011101001111111100000001110001010111000000110100010001000100010001010100010101011111010101110001001111110101010000010001001101000001110111011101000001110001000101110111010101110111110001010000111100001111110100010111000011111101001111110101000100001111000101000101110001000100110101111101000101001111011100010100000001110011110100110000000101000111000000011100110101000000010011010000111101001111010011010001010011011100110111000000000101110100001101000011,512'b11111100010100011111001111000011110100001100001101000011000001110101110000010111000011001101001101010101111111001101110101010000000011001101001100001100111101111100010011110011010101010101001111110101011111010100110011010000000001001111110001000011110100110100111111001100001101000111000111011100110100110111110000001101010011111100000011011101011101010001111100110100001111000000001111111100010100000100000011110000011100111101111101110000010101001111000101010100000011001100110000001101001111001100000011110100,512'b11011101001101010001000101000100001101110000001111110000001100000100010000010011000000011100000111110011111111001100010011000111000011010000010000000000001100001100001111001101010000110011010100110101011101010111110100010000111101010011000000000000010111010000010100010001010100000100001101000100111101000000111101110111000011111111011111110111111101110001010101010111010000001100000001011101110101000011110111001100010001110000000000010011111101111101110011000000111101011101111100011100010011110100011111110101,512'b00000000110011000101001101001101110100000101010111111111110100110000110000011111111111000000000011010111010101111100000001000111110101000100000111000001001111000100000111010101010000010011011101000100001101000011001100110100000000000100001111001100000001011100000011000011110100010111000000000101110111111111001100000011111101110101111111001101011101111101000100001111110001110101001101110011010101010000011101011101111111001100001111110100000100010001110100000101111101110001011100001101000001111111000001110101,512'b11010101010001110101110100110001110000000111010111000001010000001100110000111100001101110101010111010101001101000001010001000011110101111100110011110101010011110101001101010011110101010111110111000011010011011101000000000001111101000000000011000011010001000001110111000000011111001101110000111111010101010001000101001111010101010101011111000100010111010011000011010100000100010100001100000000010001010101110101010101010001000000110000010111010000011100010011000000010100010001000100011101000001010001010111000000,512'b11111100000101000000011100010100000100010111011100010011111100111100000100010000110100000100011111111100011101001101000000000000000000010101000100110100110000111100110111000000010111010111001100000111000001110111000100010000000011000100011100110111010000111111110001000000010000011111011111110000001101011111010011111101111100001100000100001100001100001100110000001100111100000101000101110101110000110111110100110001111100010001010011000001000101001100010100000111011111000100111100000101001111110001001100110100,512'b00001101001100011100010111011100110101000101000000010111001100000101110111110001110000010001011100010000110001011111000000000011110100111111000101000011001101000011110011110111011100001111000000010001110100011101010000000000000000111100010100010000000000000001001111010101001101110011111100110101010000110111000001110000000100001101001101011101110100111101011100000101010001010000010101010101010100110000000000010100000101110000010101000011011101001101110000011111000100000100111111111100010100000001110011110011,512'b11000111011100000011011101000111110011000001011101000011000001010101110101000100010000011111000000010111110011111101110100111100010001001100010001110101111100010011110100010001110011110011000000001100010100000000010000000111110100010111000001010001010100011100111111010100000000001111010001010000111100111100111101010001000100000100010111000001110111110000110101011101110101000100001100110101011101111100110111000001110000111111000001111111110001001111000011011111011111010101010001110001000101110101000000010111,512'b01000000011101000111110101110000010001010000011100001100000000010000110001110101111100010111010111011101110000001101000011010101011111110101001101000100000111110001110011010000011111111101010000010011000111000100110100011101010111110100010000111111011101010101001100110011010101001100010011000101000000010011010100010011110000110100110000000001000011001101000011010000110001011101010001110001111111001101001111010011010100110011110011001100011100110101001100111111000011010100000011111100000011000011110100000100,512'b00011111010011000111011100001100010011000011000000001111011111110011000111110000011100010101110111010011000000010001000011000011010011000011000100110101110001110000111100111100010011010001000001110011011100110101010011110101011100111101011111010000011111000001000011110001000000000001110111010001010001000011111100000000010100110100000101010100000101110011000101111101000111110011000000000011010011011111011100110111001101111101001101000101001111110011110000000101011111000000011111000000000101111100010101010011,512'b00110000110111110101111101000100000001000101010001000100000011011101110000110111010100111111111111010001000000010000010011010101011100011101000001000100001101110000110011110011010000110001010111110001110100010000110111001111000011110100110100010101001101011111011101011100110111011111110011011100010100000100000001001111010100110111000101000100011101001111110101000101111101000011110100011100011101000111010000011101001100111100010100000011010000110011010101110000001111000000001111011101010000000111000001000001,512'b00010111011100010011010011000111010100110100000101001111010001010000010000110001110111010111111100110000110001011111111100110011111111010001110000111100111111010111010111011100010001000000000001110101010001000011001101011111000101001100011100000000000111001111010001010100110100010000000111010011000001110000010001110001111111000011000111111101000000001111111101001100010100110101000101011101010000111111011100010101000100000100011101000111110111010111001111000100001101000101110100110000010000000000111111000000,512'b01010100010000110001000001000101110011010111110011011101110111000101010101000011010011010001010101000011000111110100001101010111010111010000010000010101000011001100110101011100110111110011110000001111110001000001111111000011000011110000110011011100001100110000010000000011000000111111000011010000000101010100010101000100000011000000000000010011011100000100110001110011110000000011110011010101000000000101111100010000011111111101001101001111011111000101001111010000000101011101000111000001110011000001010011111101,512'b00001100110000000100000000000111000111111100010000111111110001000101000101000000010011010100111101110101010011010011001101111100010001001111001101010001011111001111001101110100000100111100001101010100011101010100111111111101000011010101001101111100010111010111010011000001110101110000010000000100110000010111001100111101001111011100000000001101000101010100000011010011000100110001111101000100010001110011010011000111000101011100000111000100000000110011111111000000000100000011010101011101001111000001011100000101,512'b00110100000001000001110101110111000001010011110001000000001100001100010011000101000111010101000000000011000000010011010111000100110101000111111111000000010011110000111100001111001101010100011101000100000100110111000000000000000111010101000011010001001100111101000101110100011101111100001111010101001101010100111111010100001111001111000000010011000001000111110111010011011101010001010111010000000111001100000011011101011101010000000001110011000000001100000011110001000001011111110001011100000001001100010011000001,512'b11000001110100110001111100010101110001000000001100110101111100000001011111000000110111000100111111111111000001010111011101011100000000011100001111110000110111010100110111010111110111110011011100110101000000001111000000010100001101111100110000011101001111000001110101010001010111001100010111110000000000000011010001111101110011000111110001000101011101010100011100110101010100110101010001000101001100010100010000110000011101000111110000010111010001010111000000011101000000010001111100110111010111000100000111010011,512'b01111100110001010001010001110011110100011101111111110001110000001111110001000111010001000011000000001111001100000001000111010011110000000100110001000111111101110111111100001100000000000001011100111111111100000111000000000001110111010011000101010100111111111111000000010000000001010111110011110011111101000001010101000101110001000101010001000111110101001100010100000001000000011111000101001100111111110011010100000100111100110100110000000000110100110001010011110000001101000111010011000100110011011100110011000011,512'b01000011000100000000110001001100010100110001000100111101000011110011000001010000110111000100000000011100110101001101011111110001110011110001111111011100111100110100111100110100110000000100110001000000010000010000001100000101000100000000010001110100001101001100110100000011001101110001010111010001000001111100000011000011011101010000010011000100000100111101110111011111001101111100110001001100110000000000000111010000000100001100001111111111111111011111000001110100000011110011111111010011001100000000000000000101,512'b00010011000100010000010011000100111111110111110111000100011101001100011111110000000101010011000001000100010100110100010101010001110001000001010000010011001100010001000101000000110000110000010111110101010100000000001101001100110111000111110101000000110111000111010100000100000001000111010011001101000101110101000101000000011101010101000000001111110001110000000000001101110001010000001111010100110000110000011101010000000101110000011101001101000100000001010100111111011111000000110101000100110000010001000011110011,512'b01010100000111011100110001010101110111010011011100011100000101111100000001001100010100000111000001110000110100011111011100110001110100000100010000111111001100110011000100011100011101110000110000000101000000010100010001111111001100011100110100111111010001000100000111001111110100010111010100000011000000110000110011010111110111110001000100110011010000001111010000010111000100000001010001000100001101110001001101010000001100111101000111111101110001001111011101000011010101000000111101110000110000010001000011010100,512'b11110100111101110011000000001111110111001100111101110011111100001101000011001100110101001111010000000100111101000001111100010000000101010001000011000001000011000100010001010000011111000001000000001100011111010001000001000100000100001111000000010100000001001101001100110101001100010001010111000001110111001101010101000011111111110011001111111111000100000000111100110001000011011100000100000001110000011101000000001101110101110001111111110111110000111100110100000001000001110111001100000000111101011111001100000011,512'b00011111011100111101110000000011111101000101010100011101111100111100000011111100001111111111010011110000000000000000110001110011111101110001110001111100110001000001010001010001010011110000010001010000001100000011111101111111000001000101111100000011000111010001110100010101000000001100110001001101011100000100111111110011110001001100000000000001010111110111111101010111000000010100000111111111010111000011010000011100110001110100110100011111000111010101111111010100110001010100011101001101010011010101000100011101,512'b01001101000000000001110100010011010100111111110011110100010000110111011111000011111100111100000001010000011101110000010011111100010001001101000001110101000101111111110100111111011111000101001111010001000011010101001101110100110100110011000011010011001100111101001111010001110011000100010111000011010100111100010100010011110100000000000111010011110000001100111111010111111100000011111101011101000000001100001100110011010011110111010000111100010101110100010000000000000000110100000101010000010011110001000000000001,512'b11000000000100110001001101001101001101110000000001001101110111110011000100111111111100110011110011000101010011000111010000001101110001010100000001110111011100001100010000000001010001010001010101000001001100010011110011000000000000110100010001111100000111010111110001111101000011000000001111111101000001110000010011001101110011001100110101110001000001000011011111110000110000000100010100010111010100000101000001010100000001000001000000110011111101000100010101000100110001010001000000001100110111111100000100000111,512'b00000001110111110101000111000111000100110100110111001111010000010000111101111111111111010100110011010011000011001101001111111100000011000101000000001111111100001101111100001101001100000000001101010011110001000000001100000000110101010100110000010001000111001111011111110100000000000011110011111100000111000001110100011111011111111101010000110000010011001101001100110000110000110000001100010000110100110000010100001100010000010100001111000011110001000111010111110001010101010100110000111100011101000000010100111111,512'b11111100001101010011010001000011110101000111110100010011110000010001110100110100011100001101110111000011011101110101000101011111000101110111010011000100110000110001010011010101010101000001110000010101110111010000110111110101111111000100110111001100000100111111110101001111110000001101110011011101110111010011010011000001110001000100011101001100110001000111000000111101111111110000000101111111000111011100110011011101000000001100111111110100000101001100010100010000110101000100010100011100110100010101010011010001,512'b00000100001111000100110101000111110100000000111111010101111100001111000000001100010100111101110101110111010101110111111101111100001100001111110100001111111111110011110000010100000001000111010100001100000111011100110000111100010100000000110011001101011100111101000000111100110101011101000000110001110100010101010000011111110111010000010100000100111100001111010111010000000101000001000011000000110000000000010011000111000000010001110001011111010101000100000001000001010000001101110001001100111111000000010000010001,512'b01010101010000010101011111011111010011000100001100001101000100010001110011000011000000000000010100110101000000111100011101000000000011010000010100010111010100000011010111001111111111000011111101110001111100110101011100011101000000000101001111110000001100001101000101110000110101010101001100111100001100000101110001010100000001000000110011000001000100001101010011010100011101111111010100001100110001000011000001110001001100010011001111001100000100110100110001110111011101111101010001000101000001110111000001000111,512'b00001101001101010111000101000001000100000001000000001100010011000000010000011101000011000001111101010000010100001101000111010100110001001111001101110000110100000001110000000000000000011101000001111100011101000001001100001100001100000011000001010000000000110001110111111111000111000100110000010000000000111100000011010100001101110101011111010001000100000000010101000100110001110101000000011101111100010001000111110111111101110000000111010111000011010011011111110100110101011101110000110001000101111111000100000111,512'b01110000110100000101110000000001001111111101111101011100000001001100110000000001110001000011001111010111110000000101001111011101010111111100001100110000000101010101111101010000111111010000000011010101110001000000111111010100011100111101000101010111001100001111000100010001110111011100011100000000010111010111011100000011110001010011011111011100010001011101110100111111010101111100110000110100110000110011000001010100011101010011010111000111110011011101110101000100001100111101010100110011001100010111010001010100,512'b01011100111101010111000000010000010111110000010011000101010011110011110011110001001111011101010111010000000100010001110000011101000011011100000000000101110011000000111101010000000000001100010011011101000001000011001100010101110011011111010000010101011101000100000000000000010000111100110101010011011100010111110111000000110101001111001100000001110100001100000100010101110011000000111111011101000100111101010000011100010000010000110001010101001100010000010011110000010000010111110001110001010101000000010111000101,512'b01001100001101010001010101011111000100110111011111111101010111000011010100010000010111000100110001111111110001000101000001111101000000001100000100001111111100010100000000111100110000010101000001010001010111111101110100111101110000011101000100110011110011110000110001010011011100110011001100011100011100010000000001111111110011000001000001000000111101110101010111010101011111001100000001111100111100111101000000001100001101110011110100000111000000110111000111010011110100110000010111000000110111110000000100010100,512'b00111101000001110011000001111100001100011101111111000000010000001111110101001101000011010011010100010001110100001100111101000001010011110011010011110001010100111111110111010100000011010001000011000111110101000000000011011100010111000011011101001100000101001101110100000100010000000001110000110001000111011101111101110100000000010001110000111111000000000101000101000011000100110111001100001101001111000011110111110001001100000001010001010111010100011100001101111111110111001100110000000001010011000111000001010001,512'b00011111111111000000000000110000001101000011010011010101001100110000110100000000000001110001110001000011110011000101000011110011000100011111010011010011000000011111110101010011010100000000001100000101001100011111110101111101011111110100000111000011010100000000110101110011000000010001010011011111011100111100110000010111000011010111110011111101111111000101000101111101110001111100111101110011000011000100010000110000001101110000010000111101001100110000111101011100010101110101110001001101110111000000000011000001,512'b00001101111111111100000000000100111111110000000011010011010011110100110101011100011101011101000101111100000100111101111101000011000000000000000111010000010101011111010101000100000011111111000001001101000101111100110001000000010011001111011111110111000000110111111101111100000101111100010011001101110111000101000011110100001100110111000100000000001111110001111100000111010001000000010011010111111101111101110000001111000101001101000000010011011111001111110000001100010100111111010001110000000101000000110001110101,512'b00110011000001000000010101000011110101010100010111010111110111001100011100001101110101110101110101000001110011111111010011001101110100001101000001011101110000111111011111011101011100001100011100110111010100010011011101110011000011010011110011000001000000011100110011000000000011011100010000000101011111001111001100110100111101000001011101111100010100001100000100010111010111000001010000000000000000010100110000001100111111000101001111011111000101000000001111001101110001110000001100110000000101000000110101111100,512'b00010101001111011111011101110101110001000100001111110000110101011100000011010100110011000100001100010001000001110000010000110000010001110101010101010000110001111111000100010100010111010001011100011100111111011111011101001111011100000101110000000111001100110101110000110000000100000001010000000100010101011111010111000100110001110100001100010000111100000100000101001100011100001100000101000101011100000111110011111100010001000001011100010100110101110001001111010100010101111101010011110111001101111111000000110100,512'b11110000000100011111110100110101110001111100000111010000010101010100001100010000010011001100110101111111110101001111000101001100010011000000000101001100010000010100001101001100111100011100000001001100111111111111001101010001110001010000111111110001001100011101111100000001000001110111110000011100111111010000011100001101000001000100000000010001111111010000110011110100001111110111001100111100010101011100110011001101011111110100000100000000011101011101001100000100110111010100010101001111000000010011011100000000,512'b01011101000111010111110111111101000001000101010000010000000011010111110000111101111100011100001111000001010100011101010111001100010011110100110101010011011100001100010100110111010111111101000000110001011100000000110100110100110111000000110000111100010101000000010101111111010101000001000011000011010111110001011111001111000011010001011111011100000111000000110000010000000100010101110001011100000011000100010000000100000111001100001111010011000000110001010111110000110000111100000100110111000001001100010101110101,512'b11000101110000000100000011110100011100010100010100001100110000010000001111110101111101001111000111001100000000111100000011010000011101000100001111000001000001000011111100000100010000001100110000010000111111001101000000010011010101111101010111010001010001000011010111010001000011110111110001000100000111000100110101010101010100110111000011010111000011001111110100110001000101001100000001110101000000001101000101000111001101011111001100000011010101000011010101000101000011000011001101011111010100111100000001010000,512'b11000100110001010101000000110001010000111101001100010001010101001111000001010000011101001111110000110101001101011101010101001100011101000001110000111111001111000111010001111100001100010001110101010000110001010001000000000011110000110011010001001101000011111101010011000011000001001111000000110000010101000101111101001101010000001101001101011101110011001111010100000101111100001100110001011100111101000011001100110101000000001111110101000001110101010011010101001111010100000111010111010101110100000101110111110000,512'b01010001000100110111000000010000111111010000000011111101110101000111010001000011000011001111000111110011001101001100001101000101011101011101010000111111110000011100111100111100110001010111111100110100011111111111111100010101000111111100000001111111000001010101010000010000001100000111000100011111001111110000000000011111110100010101000000000101000011010001010000110011110100000000010001110001001111011100000101111101010101110111111111010111000100000001001100010011001100001100001100000100000001000101110100000100,512'b11010011110100110101000000011101011100010101010001000001110001000011010000000100110000010011000011011100110011110011000111110001000100000100011100111100000000110100110011110001010011001101000001111111000001001100000111111100000111111111010100110101110000111100010001010101110011000100001101010101010001111100110101111100000111001101110011010101010001000001010000000111011100010100010100000011110001000100111101110001000101010011000100010011110000000011011111000000000111110001000001000111110101010101110001111101,512'b11000000111111010101000011110100000100010101000000110000011101010111000000011101010000110100000011000000000100000000000101011101010001000100000101000101000111111100000111000101010011000101000100000100111111111101001100110000001100001100111100111100111101000100011101010111001101010101010111110111010001110001010100011101000111011101000011010101011101000101111100000001111100000111010100110101110101111111001111010111010000000011010011110000010000011111010001110101110100000011000100010011000001110001000001001100,512'b00000100011101111101111101011111001101010111010100010100110000000001111100010011010001010100010101001100110000000000010100000000000101011100110000010011001101111101111101000111010100000000010100011100000001000000011101111100010011110001000111111111001101001100011100110100000000001100010000110011011111111100001100010100001111111111110101011111000101001111110011001111110011010100110000010011111101110001010001110100110011010001010000011111000000000101000000000100011101010101000111110001110100001100001101010000,512'b00010100001101110000001101000000110001110101010001110001111100010011011111001111010011111101111101111100110100010001110100000011001111001111010100110001011101001100000011000001000101000000010101000000000011010111010001001100111101110101001101010011110000010000001100000101011100110111001100111100010011110011111100011111000101010000000011110111010011011101010001000100000101000000011111110111010001000011001111011111000011011101011100111111011101001111111101010000011111110101000001001101000000001100111111011100,512'b11011111010100001111000000011101011100111111110011000101110100110011110100111111010011000000110101001100110100010101111101000101010100111111010101110100000100110011110100001100110100000001000111000001011101110000010111110101011101110000110011111101010111000001010001000111001100000101110000000011011100111100010011010000010101011111000101000000110001011111001100010100010100010100011100010000001111001100110100110001010100110000010100000100000011010100011100111101000011001100110011110001001100000000110100110001,512'b01000111110001110001000000001111010000000001010000011100110011010011010001000011001100000100010111011111000100000011111111010001011101011100000011000111010111001100010000110011111111000101110100000011000001011100001111111100010100000111001100000111110000011100011100001101010011111101000000000011000011000001000101001100001101110011010000110011010100000111110101111101000111110000111100110101000011000000110000010011011111000000001101011100010011000001000111000100011100010111110100111100110000000001000100000011,512'b11110100010001110011001111000000001100110111110011110111010111000011011101000111000111011101010100010000000011110001000001110101111101010111110101000111001111000111011100110000110011111111110100000101110100001111010000001111111100010011110100011111111111111111010001110000000001110101010000000011010100110000000011000101010011010001000101010111111101110001110100110111001101001100000100001101011111010000000001010001111111110000010001000000000111000011000000110111110011110000110111110100010011000000110100001100,512'b11010011000011000111011111011111000011110000001111010011000100001111001100010001110000110111010111010100000001000001010000000000111111010001110011110000010000111100011111001111000001010100000100110100110100000011110000010000010101010100110000010100000000010001000011000011110101010000000011000000000001010000011101010100011111001101000001000011000011010111110111110000000000010101011100010100010111010001011111011101011100000101001111011100111101001101000001001101010101010000001100010000010001010011001101010100,512'b01000011010001011111000001110011000011001101001101000011010011001100110111010000000101010000010001000101010111000101000101010011011100000101010000000101000100111100000011110101001111010011001101011100011100000000111100010111110101110101111101010101001100011101010100110111010001011100000100000001010101011100010001010000011111111101000111011100011101110001001101001101010000011100010111000101010111001101000011000011010001000111001111111101000011110100010000010011010000110000110001010111000100010111111101000000,512'b01010100010001001101011111010101001100110011000000110000010011000111000101010101011101010000010111001111010001110001010100110001000100110000001111000000010111110000010011000100110000110100111111000001010001000011000111110001010111110101000001011101001100010000010111010100111101000011010011110001000001010111010011000000111101010000110001000001110001110011011100010011110001011101001111110101000000000101010000000101010100000001001100110000000111001100000000110011111101110101111111000000000000010000111101010000,512'b01010000001100000111011111010000110000011111110001010001001101111100000000010000010011110101111101010011000000110100000100110000000000110000001101000000001100000000110000110100000000000011110111010101110100111111010100110101110011010000110001000001010000000100110101110100110000110011001111001100010000010000011100010100111101000101010101011100000111111111000000110100001100000000110000010011010011010111010000110001011111000011110001011100010011111111010011011111000100110100110011011100001100110101000101010000,512'b01110101110000011101110101110100110011110011111100001100001100010100000111011111000001010101011101010000111100000100001100110011000000000111110000110000011100011111010011000111111111111101010111001101011111000100011101000000000001011100011101110011000100000001110000000000011101000001011101010000011100001100000111110100010101001111011111000001001111000011010001010100011111010001110101110001110011001101111100010000010000111100111111001100111101001100111111010001010011000001111101010101010000111111010000011101,512'b00000100011101000100111100000000000100000000011101010011000100110101110000010011000101010011000000000101111100000111010011000011110100001101000100000000110001000100000001011100000100110011011101000101000101110111110011001101010001110100010101000000001111000001110011000000010001110000000000010000110100111100010100000001110111110001110111111100010011111101001101110000111101000111000111011111010100000101000101001111010000000000010001010111011101110011010011110000010000011100011101000000011100000011111100110100,512'b00010000110101110001111111000001110000110101011111010100000000010100000001110011011101000011110000000001001111110101000000111111001100011111001111010000111111010100110100001101000100110111000011111100000111010011000011001101000000110111011100110000000101110000110101011100000111110000000001010001011100000011000100000011010100000000000000010100000100001101010111110111111111010111000011010111010000010000000111111100000111001111001101000101010011000111110111001101000100010001110101010001011100000011110111010000,512'b11011101010011111111010111010000110011000011111100111101000101000001110011000111110001000000000011010000000000111101110000000001010111000100000111010011010100001111010101010011110001011111110100000100000001010100111111011111000100110000110011011100011111010000010011110000010011110101110000011111001100000101110100001100001100110101010001110101010100010100000000111100000011111100110000111101011100010100011111010000110111010111001111011111110101000011000000010100011100011101000100110111000000001100110001011100,512'b11000000001101010000001100001101000001000001110000110101110011111100010001000101000001000001000111000100111100010100000100010101010011001100000101110000110111000101001100000011010001110100000000110111110001000101111100111111111100000100011100000011001100110011001101000100000111001101000100001101001101010000011100010100111101011111110100000011000111000100000111110100000001110011000001011101110000111100001111000100110000010100110000111111010100011101000001000011001100000101010111110111000000011100010111000001,512'b01000100010000001101000101110001010001000100010000010000001111001101000100110000000111110101001101110001001100110111001101010001010001001111001101000111010101001101111100110101011100110011001100111100000111110100010100000000001111000001010101010111010000000101111111010011110100001100011100011100111100010111001100110111001101111101000000110000111101011100000100010111110001011111011101010100000001011100110111010111000000111111001101110101111100010000110100110111010101111101000101000100010011010101000011001100,512'b11010000000011000000010111000000110000000100001111011111000000110101000001010001001111010011110100010000000100111100011101011100110011010100010111110000010000001111010101010001000001010000010001110100011111010111000001010000000011000100010101010111000100001101000011111111010000001101000101110100000100111100001100011100000000111100010100010001111111000101111100001111000000001100001100110001000111111101110111110001010111000000010001110001110100000001110111010001010101000100011100010001000100000100111101000011,512'b11110100010011001100000001111100000011010100110111011100010011010011110001110000001111110111111111110100010100001100110000110111010101000101000111001100110101110001110111010111000100110011111101000111000000000101111111010101011100110111000101010101110100110100010111011111000001110000110011010011110000110111110000110001110011110101111100111111010111010100000000111111110000001101111101110011001100110111001100000000110100111111010100110101110001010111000000010001011101011100000101000001010000110111000001001100,512'b00001101000100111111000000000001000111000000000001010001110111011111001100000000010000110011110100000001010011010000111100110000010000110101000001010100001101010100111100010100011100110001000100000100010111000000111100000100110011110111001101111100010001010001111100010100000000010000110011110001010000010011011111110100000100110001111100001111000000110001010111010000111100011101011111000101011100010000000101000011000001110000011111111100000100010011000101010100001100110111000000010001010100000000000100010100,512'b11110000110011010001011111001101000001001100001101010001111111010000001111110111000011011101111111001111000100011100000011110001111111110100111101010000000001011111000011011101010001010000110100000001111100110011001100110011000111000111000111001111110000010111000011010111010011010001010100010001001101010101010101010011110000110001000001000100011111000100011101001101110100000011010000000100010111000111000000000111010000000011110000110011011111111101000101011101111111010000000111000100010001000000110001010000,512'b00111100000100110101000000000000010011001100010111011100010011110100001100000011110000000100010011111100110011010011010011000100011111001111110111110111111100000001000001011111001101111101000100010101001100001100010111001101010000110000001100000001011111000011010000001111110011000000000100000011110100000100011111110011000100010101001111110011111111110101110000000101000100110111110011110111110011000001110001000011011111010001000101000100000111000001010101010011000001000001111100110100010001111101110011111100,512'b01010111110000000001000011011111000001000101000100110011011111011101000011110000001100111100010000011100000100110011000011111111010011110001000011000100000000000101010001010000011101001100000111110101110011000011111101001100110001110000010101001101011100000100010100010001000011011100000011010011111111010011010011001100010101111101010011010001001100011111001101011111011100001100001101001111110000110100110011011111110011010011000000111111111111000001110011110000111101000101010000110000000100000100011111010111,512'b11110111011111010100111111110011000100110100010000011111000111110111000001111111000001110000111100000100000001001111110000011101000101010000010000000000010100110111110100011101111101000011110001000101010100001100001111000101010011011100110101000111010100000001000101110000000000011111010000000100110101000001000001010111001100111100110011011100001100001111110111000100001101001111000111111100000111011100000100000001010011010001010100001111010011010000110100000101110111011111011100010101000011110001111100010100,512'b01110100010101010000110000001100000101010000010001111100010100111111011101110011000111000100010011000101110001110111010000010001110100010111010000011100110111010000000001000000110001001111110100001100110111000011000100011100001101111101010011011111011100010101001100010000010011001100000100010011000101001111011100000100010000000101001100010111000101000000111111010101110001001100011101111100010011000000010100000100001100110011001101110011011101010101000100001100000111001111110000110101000000010011010111010111,512'b01001100110011010001000011000100000001000001000100000000000011011101111100010111000111001111010001110101001101110101001101010000000101000011110001010101110000001111110101000000001111000001000100011101110100000001001100110001000001111101110000000101000000000011011101110000111101111100011111001111110001111101000001110011110111011100011101011101010000011111110000001111110100011100011101010001111101001101111100000011010011110001010001010111111111111111000101000111011101010101010001001111111101110011110001110001,512'b11011101111111111100110111111111010001000000001111010011000000000000110000000100111101001101000101010111010100110000110101110011110000011100001101000000000100110001001111010001111100111111010111000101000001110001010101111111000100110000011111000011010000011101010111001101010111000000110100000100000011010011011101000100110101001101000001010101010111111101011100010001000001011100010011000001010101110100110101001100010000011100010011010100001111010100111101010001010100001101010101000000000011010000010100110011,512'b01010101010100000000010101111100110001000101110000010100000100001111000001010011011100010001001101011111011101010000110101110000010100010000000001000011000011110101111100110101110100000011110001011101110100110100111100110011001101000000011101000111010001000000000011110000010001111101001100111111000101010111110001110101110011111100000000110001011100110001110100000101111100010011110111110100110101110100010000001100110001010011000011000001110000010001110100001111001100000011000011000001000011000011000111110001,512'b01010111111111000011111111110000000000010011110100010100001101000001000100000100000111111111011100001100010011000100001111001100000000111100000011000000110100001101010011000111000001001101001100010011110000110101011100000000010001000111000011001101110111010000000000001101010111001111001100001100010000000100111100110100011100010000010100000111110101110101000011000001000001110111000001001100000101110011010111001111010100111101010011110101010101000000011111010000000011010101010100011111010100000011011111110000,512'b01111111011101000001111100000011110000110101111101001100011111110101000101111100010000010100001101110000110000110001110000010111000000010100000011000000001101011111010000111100001100000001000000110000010011000111010001001100000101010100111100110111000001110101000101010100010111110001010001000101111111010001010011110101011101000100111100111100000000000011001100011100010111010101000101000100110000000001010100010100111100000111001101110100011101011100001100110100010000001111000101010100000111011101000011010100,512'b00010011010111111101000000111101000001001100010011010000010011110100011100000111110001110101000111000101110100010000010011000000010000000001000011011111000000001111110111000001000100010001010100000101110001110001110000010100010101000001010001110001011101001111000000001111010000000101000000010100111111010000110000000100001100000100110101000011000000010011110000001101010000110101000000010001110000110011110101110111110001110011001101110111110111000111110111001100001101000111000101010011010100110111000111110100,512'b11000111000001011100000000110001011100010100110011000000110011010011010011000000010011111111111101000100111100010101110100011100110101110001111100001100110100001101000000010101010100001100000111110011000011110000001100010011110001001100110000010101010101111101001101001100001111001111010011011100111111000100010111011101010000010111000111011100010000010101010111000100111100000000111111001111011100110100110100011100011100011101000000000111010000000111110101010011000011000001110001000111110001110101000001110100,512'b01110001011100111111011100111111000011010011110001000101000101000000110000011101000100011100000101000001000001110011110000010111110111111100000000010100110111010011000000111111010111110111010011110101010100001101110011110000010101010111111101000111011100011100010101010011000011000100110100111101111100110000001101001101010101011100000001010101010000010000000111000000011111010000010000001100010101001111010111010101010101000000010011000011111101010011000101000100000101011100011101010101110100001100000101000100,512'b00010111000101111101010011110000111101111100111111011111111111000100010101000011011100000111110011111100111111011100000001010001000011110100000001000101001100110100111101000011110001000011010000001111110111110001110000010001011100000100010001000011010111000101000000000100010011001100000111000000110000010101001100001111011100010000010000001101000001110011110000010101110001000101001100000000001101000011111100010100000101000000000011010101110001000000010000000011001111010100000000111111010011111100110111000001,512'b01000001001111000011010101011100110001001100000100111100000100000100011100110000001111111100001111110100000101010001110111110011000000000101110100000111000011010000000000111111000100000101010011000000011100001101001100110001000100010001110111110000011100010011010000011111011111110011001100111100110000000011110001110100000000011100000101111101001111000011110101000000110000001100111101010111110100110111000101110101010001000111010101010001001101000101001101010111011111111100111100000101001111000011000101000011,512'b11110100001111001111001100000100000000000011110101011100111100111101111100001100010101000011010011011101000011010001010011010001010100000001110111000011111111111111001111001100110000110001110001111101110100111100001101000111001101000001000101000100110001110011001100000100010111000000110100011100110100001101000000000111001101110011000001110111110000111100111100111100000000011101010000010101110000010001110000010101010001010000001101110111110011110000010100110111011101110001010100010001000001000111000011001100,512'b00000101010101010000010011000000010011000100010011010100000011000101111101110011110000011100111100000000010111011100010001110100110111010000110101111100000100111100010000000000000000110100000111110000111100000101010000110011000111111100110111010101010100001100000111001100110100000000001100110001000111000101010000110011000100010011010001000000010000000100011101110011110001111100111100111111000000000001011111000100011101010011011100001100000100110000010001011101000111000100010001111101001100111100010011000000,512'b00110000110000010011011111001101110100000000110001000001110001010111000000011101010011010001011101001100000111010111011101111101010011011101011100000000001101000011010111000000000101110111010111110001011101110001110000011101010100110001001111011100111111110001111100010100010000110000110001110011111111110000001111010011010001000100111100110001110000010101110111110100011111010000000000000000111100000100000101000100011100110000001101011111001111000011010100111111000100000100000111111100010101111100010001010100,512'b01000011011111110000001101110101010000111101010111110101110011111101111100011111010000010000001101011111110001000001110011000000000000010101001111001111001111000001001101000011110011010101000011000111001111111100000001010111011100010011001100001100000000000001110100111101111100111100111100000100110111010011000000110111000111110001001101001100011111110011010100000001110001000101001101011100011111110000011111001111000001000001010011010001110001011100001101110001110101001101001101011100010011000111011100111111,512'b00011101010111000000111111110000001100110100010111000100000011000000001111010011001100111100000111000101000101000000011111001100000101000000111101110101110100010101010000110100010000000011001100000100001111000111110101110000001100110001000000000001010011000000110101010000111100001100010111110011010001000100111100110001111111010101000101000011010011001100010100000000010100000011110000011100000000001101000111000101000001110000010011010111000000110100001100001100000101010011110011110011010000110001000000110101,512'b01010001001101111101001101001100000001110011110100001111000011110100000101010101110000000111001100011111110100001111000101000001010011010101110001001111001100110000111101010101011101000001001100110111111101010001000001010100110111010100110011010101000111111101000001001101001111110011111100110100000000010000111100011101111100010100110100110111110101111100000101111111110101000011110000000001011101110100001111001100110101110100111100010100001101110011110100010100010101001101001101010111011100011111110101110000,512'b01000000011111011100010111010001110001000000001101111101110011010011010100000000001100010000011111110000111111000000000101110000110000010000010001000101001100010101000101000011010001010001110011000001000000111111000101011101000101000011111111000011110101000001011111010100011111010100000100111111000000110011110000000011010001110001000001010101110001000100000101000100110100010100001101000011010011110100011111001101110000110100000011000011010000010111000001111101000001001100001101110000010111011100110100000101,512'b01110111011100010000011111000000000100010101011101000111010111000111110001001111110001000101000011000000010101111101000101000011010111110100110100000100110111001111110111001100010100111100000111110100111111001101000100010001000011110000110001011111000001001101000100110001000001110101010001000101110011010100111101110011000111010001011111110001011101110100011101001101010011110000110011010001110000000001111101010001011101011101000001111100110011010100001100111101111101000100000101010100110000110100010011000111,512'b01010011001100001100110001000000111111110001001100110001110111010001110000001100001111011101110001001101110000011111110101010111111100000100110011110001011101001101011100111111010000000100001100010011111101010111111101011101000001010000010001110100010011111101110101110101000011110001001100111101000100111100000101000101110100000101111101111101000111010100110011110000001100000100110001110000011111110111110000010000111101111101011100000101110011110011000001000000001100010100110011111101110001110111001101110001,512'b11001101000011010111011111110000110000010011001111000011000000110111001100001111011111011101010111110000001101001101010000001100000101000100111111111111010111000011110100000100001101000000111100000101111100000000001111010001111100001101000000011101111100000001000111110100111101000101000111000001110100001111111111110000011111010000000001000100111101011101010000011100000100110011000001110000000111000100001100010000110001010011111100011101000111110001000101110001111100010001110011001101010100000011110011111101,512'b11011111111111000000010111000001010101000101010101110100000101010101010000110101001101000100000100000101010011010011110111011101001100110100010011000101001111000001001101000100011101110011001100110001011100110111110101011111010011011100110000111101110100011111010000010011111100000000010011010100000100110101110111001101111100010011010000110000111100010100011100000011010000000000010101010100011111010001010000110100010011110111111100001111000000000000010000011111010001110100110000110100110100110100000101110101,512'b11000001110011000000110100001100001100000101001111000100000100010100010100000111000100010001110111001100011100010001110101110100000000110001011100001100000111000011010101000001110101001111010101110001000001010100001101011100110001000001001111010100110100000000111101000000000000001100010001110000000001000111011100110011011111010011110111010111011101110101110100110001010001010011011100001100110001000101010101000011111100011111011101111101010001110111011100001111010111010100000011111101000101011100111101000101,512'b00000001000001000011111111000001000001001101000001000011001100000001011101000011010000011101110000110001110101010011000000001100111111110000011111000011010011011111010001011111011101111100000111000011000101001100110001010000110011000111000001000100111101010101010100110000110011001101000111110111010011000100111101000011001100000101000000001100001111011111110001110101010101110011000011001101000100110000000000001111010100000000110000010011010100011100001101001100011101111100110100000011010111111100110011011100,512'b00011111110011110101001111110101001100010001010111110111001100110001110100010001110001000111000001110001000001110101111100110011000100001101111101010100000001000101010011010011011100000001110000000101000001011101010000010111110111000100000000000100001111010000010000000000110101011101110100000011000011110100001111010001110011000100010011010100000001111100000001001101110100000100110111000111010001010011110100000001001100110101001101010001000011111100010001010001001101010101001101110101000001011111011100001111,512'b01111101000101110100000101111111001100001100010101000101000111111111111101110111001111011100000011001101110001000001000111000111110001000100011111010000110111001111011100111100010101010011011100111101110000110011001100000011111100011100010100011101001100111100010101001101010111110000010011011100011101000001001100001111011100011101000111110001001101001100010101110111000000000011011111010101110100010100111100001101000000000101000100000100010111010100010011000000111101111101011100010101010111000101011100010100,512'b11000001000100110100110011000111000001000001000000110000010000000000001100111111010000010000010100000000110100011111111100000101010101001100000000010100001101010011000000110000011101000100000111110011110000111101000111110001010011000011000111110111000100001111001100110000010111000000011101010101111100110100000100000001010100111100000011000001000001111111000111001100000001001100010111000101001100000011111100000000111101110001110001110100000101010001000111010011000011010111001111110111110000111100011100110001,512'b11000000000011000011010011000000000111011111110101011111001101010011110111010100010100001100110001000000001100010011010100110011010111000101010101000100000000000001110101110011010011010111010101000000001111110111001100000000010100110000000011001100000000010011011100000100010111111111110111110000000111001111010011000001110100001100110111110000011111010111000011111111001100110111001100011111110000111101110101000100010000000101110001010001001111000111011111001101110100010101000000011101000100001100000101111101,512'b00000111110001011101111100010000000111010101000011110101111100110111001101001111000101010001001100000111000001000001011100001100000011000101110000111101011100110101110100110100010000000100010000000011001100000000011111110001110001001111010111110000010000000111110101110101110011010011010000001111001111000100110111010111110100000111011101001100010100000111000111010011111111000100110000000100010000111100010100110100010001011101010011110000110100110000000100001101001101000011000011000000000101110100110000010011,512'b01110000001100110101011111000001000011010000111100110111001101000000010100001111010100110000001101111111000101000000000000110100000111011100000100001101110100001101000111001101110111010100000000000111110000011100011111000100000100001100001101011111011100001100000111110001010101000111000111000001110101001100110101010000111101001101110100010100011111111111000011110111010011001111011100111100010000010101010100110111001100010101011101000011111100011100010101110011010100000011010101110000110101010000010011111111,512'b11011100010100010000010111111100111100111101011100010000110100011101110100111100111111010001110001110101000111001111010111000101000000001101110000000111000101111100000100000100110001000001010011111100000011010000010101010001111111111101111111001100011111001100000011010011001111000001000001110001011101001100110000010000110100010000111100010111110101001111010111111101001100000011110101000011010001000111000000011100000111000001110000010000110001110101010001111101010111011100110011011101011111000000001100011101,512'b01000000111100010000010111110111111111000100110111000111111100010001000111001100000101110011001101000000010100001100000100001100010001010101010000000011001100111101110001111100001111110100000001010001000111000011110100011100110011110100110011010000000000110101111101010100000111110001010111010101001101011100000100110001001100000001001111000000010011000111000011000001001101001111110011111100011101010000000100001111110000010100110100010000000101011101110111110101000101001111110100001101110011000101001111110100,512'b01000001001100011111001100110100010011110001110101000001001100000001000111000111110000110001110100110011111101001101010100001101001101000001000000000111000101110011000001110011000100010011001100001101111111010000010001010000001100011100110011000000010001001101000001011100110001110011110111000111011111010101011100110000001101000000110000111100001101010111001100001100000101000101010011011100000101000111000011111101111111001101001100001101000100000100000001000001011111000100000111001111000011000000000111001101,512'b00000011000011010011000101000001011100011101000001011100010100000111110000110011110100010011011101000111000111000101010101110000000111111111111100000101000000110101000111000001011101010101000111001100110100000011010011110001111100011111000101000101000111000101001100000111000011110001010000110001000111001111001111110100000011010100000101110101000000000100000001000101110001010101000000000000010000110001010101000000000101111101011111110111111101010011110011001100010011000000110111110001010111010001110111000101,512'b11010000110111000101010001110111110101000111001100011100000111110000000001000100010111110111110100010011000101110100110000000000001111011100110000010111000101010001000100001100010101111100000100000101001101011100000101010100000111110001011100010100010011010000010101111101010000000000011111000000000000000100000001010111110101000001000001001100000001010101011111011100000000010100111111110011000000010011010101001111000111011101111111001111010000001100000001110000110011001101000000001111011100110100000100011100,512'b00010100000000111101010001010101000011001111010101111101000000111100000011000000000011110011110111000011000000010001010000110111000001110011011111110100111100110111011101010100010111010100010001000000000100000001110100010111010000011100011100010000000100010011010000001100111100010001001111110001111100000001011101110100110000011100110100010000011111000001011101110001110100010111010100000000111100110101011101010011000101010111000000000001110100001100110101010100001101000101001101010000011101010011010001000011,512'b11011111000001010001010000010100110011000011110111110011001100010101000100110001000111000011011101010100011100011101000011111111111100000101110001000100000101000011110111000000010111001111001101010000000001010101011101110111110100111111110000110100000000110011010011010011010000000000111100110001010011011100010000001101010111011111000011000001010001000100010111000100010000111101000100010011010000110001010000010101110111110100110000000000010011110101010001010111000011010001110000110000000100010011001101110011,512'b00110000001101111100110100010000110111000001000000010100110111010101111101001100001100110000111100011101000111110001011111010101000011111111110101011111010011000011000001001101010001010000111111111101000011011100000000010111011111011111000101110000110111010100110011000111011101000000111111111101110011000001011100000011110001111111000000010000011101000000000000000100010100110101000111001100000001010001000111010100010101000111110100111101010000110001000001110011001101010100000001010111000111000101010100001111,512'b11110101011101000011111101010100010001111100110001000011011101001100000011010100000101000101000000000011111101000001010011010111011100110101011100001100010111001101110111011111111101001100010100011100000011000011110000010111001111000000110011001100000000010000000100011100010100111111011111110000000011111101000001111100000100111100111100000001000000111100001111011100110011001100011111000011000100000101000111010000001111000100110011000000000011001100000011110001001100110011000100010101011100110011000001000011,512'b00111100011111110001000101110111000011000011000001110000011101001101000000111101011111111111010100000000000100110100010101000101011111010001110101111101011100001111010001110000110011010100010000010111000001000111010111111111000100010000000101010001111101010111010001110100010001111100111111000011110100011111000101000101000001110000011100001111010001010111111100010001110011001101111100011100001100000000011100011111010111011111001101111111110011000111110101000011011111001111110001000100000011110101000001000001,512'b11011100000000110000111101011100111101111101000001010111010011001100000001000011111101000100011111000011011100110111000111011100000011000100110100000001000111000111001100110111010011000101011111000101110001010111011111010111010011110100010001000001111100011111000001000000010001001100011101110000110100010100001100110000111100000001111100000000010000000000000100001101110111111100110000010000010001010100010011000101010011000011110000010001000100010100000011010100111100001111001101001101111100010000010000011100,512'b01011101010100110011000001000011001111110000110011001100001111000101010111010011001101000100111101000000000000110101111101010101111111110000011100000111001111110011110101110100110001000001001101001111111101010011010000000101000111010111000101000000110111010100111101010000001111010000010100110011011100000111010000010011010100001111000111001100000000000001110100111101001111010011111100111101011111011100111100000001010001010001001100000001111100110000110100011111010000000011010101011111011100110111111100010101,512'b00011101000011001111110100110101001111011101001101110000001101110111010000000011110100011101110100010011011101000100000000000100110011111101110100010011001101000011001101001111010100111111010111110000110111000111001100011101000001010000001111000011110001110100001100010100000001001111000100111101110001010000000000000001000000010001001101001100010111001101000000010100000001110011000011000011110001011100000101001100110100000101000101000101010011000111011111010011001101111100000000001100000100010011000111010001,512'b00000011010000000011001101010000110100010100001100111111000011110011000001000011110111000001110011000101111100111100000101000111110100011100110011110101000001001101000011111101110001000000011111111100000001000100111100011111110000000000000001110100011111110100000001000011001100000000011111110101011111001100011100001100111100010001001100010001110111110000001111110101000000110100011100110100000111001100001101000000111101010111110111000101110000010011011111010011110000110001000111000001001111001101000000000000,512'b00001111110000110100110000111111010011000000000011111111000100111101001100110100000111000000010001001101010100011101010100000100110111010111000011010011110001000101001101000000010101110001000111010001010001001101110100000001110011000101010000000000000001000100010011010000111101001101011111111100010111110001110101000001110111111100010000010011010100110101000101001100001100110101000011000101111111001111001111000001000100110011001100010101110111110111010100000011011111000101000111000000010011010111000111111111,512'b00010000110011000001000101111111011100000011010001010000000000010001000000111101010100110011000000000111010100010000001100110111001100010100001111000011010101001100011100010101000001110101110100001100110000110001000011000011000001110101110100010100001111010001110100010101001101110100010011010011111100010111110001001100111100011100011111110011000000010111010000110000000001010101010001110100011111000001110111000011001100010000000000010011010001011101010111111111000101110000000000011111110000000111010100010000,512'b01110111000011110011010100011100001101110000011100011101110011000100010000111101010001110001000100000001010001110000000011000000110100110011010000111100000111110000001100011100111101110100000101111101001100110001011111110100001101000001010000000001010011000101110011010001010000110000010111001100010100110001000000001100010011111100010101111111111101000111110111110000111111110000001100110001001111111111000101000011001100011101000001001101010000000000111100111101111111000111000011111101011100010000111101011111,512'b00010011011101011100000101011100000000011100110001001100011111001101000000111111010000000111110100010101000111011100001101011111001111110000110101001100000100110001110101001101111100010001000101010101001101110000001111000100110100011101001111010101010101001101001101010001000101111111000101001111110011111111000000000000010101000000000001110011000100000111010000111111011111111100010011111100110001111100010000110101010100010100011100000101000011010001000000001100010001000101010100110111010111010100001100110001,512'b01010000001111000000110000000011010001000001001111111100001100000011001111000001110101000101000000111111110000001100000000011101110000110111000001110100010000000011110111110101010101000000000000001101010001111101110011001111110100011100000001110011010101111100000011111111110100001100001100110111110000000011011111110111000101010001000001001101110101110111110001001111110111000011010000111100000100000111110101011100110011001111110011110000001100010011010111110001000011011100001100110100011101010000000001010101,512'b11000000111101110011000101011101000101001111111100110011000111110001110111011101111100110101000101110100010101011111001101001100000001010101110001000000110000000000111111000011010011000011011100000011000101110011010011010100000111000111010100110000110101011101001111111100010101000000000111000000001100110000010100111101000100110001001100111100111100010001111101001101001111111101000000010011000000000011000001110011000100111100011101001100000011010011110100010000110101011100110100000111010001011111110100000111,512'b01010111000111010000010000010001010100110000110100011100000011000101010100010001010011111111110101011111110000110101011100000011000111110111110001111111011101000100110101110011000100010000010000010011110000000001110111000011000001110111010111000000010011111100001100111101011111110001011101010000001100000101010100110011000000001111001111111101010001010111010001110000111111001100010000010011111101010100110001001111110011001100010000010101000000111100010111110100001100111111001100110000110111001111110000010000,512'b00000000000000011100010101110011010101110001010001110001000000000101001100000100010011011100110011001101001111010001000101110001110000110100001111010101110011010111000001111111011101010011011100110001010011011101001111111100001101011111110011010000110000001100111100110100000011110111000100000000000001001100110111010001111100110000001101000001000011110000001101011101010000110111110000010011110011111100011100001111001100010000111101110100001111110011011101001111010011110100000011011100110011110001110111001111,512'b11010100110000010001110000001100111101011111111100010101001100110000000101000000010001010100010101000011011100000100001111000001110001001111010000110001001100011111111111000000010000000100001100001111010111110111110111000100001111001101010100010011001100111100000111011101111101111111011100010000011100010011001111010111110011010100010111111101011101010101000011010100010001001111000001110111000000111101000001111101000001110011001101001100111100010001110000010001110001000001111100000011000000000100010100000001,512'b00110011001111110011110100000000010000010101000100001100011100000011000101010001010000001101001101000101111100001101000111010011001101000011011100110011010000001100010111010001000111110011001100010101001100000001000111110000000000010011000000010101001100110101000001001101010111000100010011111101001111110011110000000100110101000100000100111101010011110011001100000001011111111101000011000001010101010100000000010011000100001101110011010100010100010000000100001101010111011100010011001100110111111101110101000011,512'b01011100000001010101000000001100111111000100011100110000010100010000000111000100011100110111011100111100000011110111010111000011001111110001010111110101111101111100011101011100110011001111011100001111111111110011111101010001000011000000010101000011001101010011010101001101111111110000001111001101000000110000011111110011000011110001010100000111110100110011110000111111110001010011110101000111001100000100110001110111001100010000000000011101110001110100111111010001000101110100010000010101000000111111111100000001,512'b01010000001101000000110101010100000001010100001100110011000111110011001101001111111100110111010111000001110011011101110100010101001101011100011111110111011100011111110111111100000011010100000100010111111100000000010001011101000101000001010001010001000111110011001100000011000000000000000011011101000011001100110011011100010101110101110111001101001100010111000011110001000001011100110101000001010101000101001100111100110000010111000011000011010100000101000011110101110111110111110001000000110101111100000011111100,512'b00000000000101011100000001000101111100001100110001000000000100011101000000111100010101110001000011001101010011001101010000010000000011110011000000110100111101010100110101000001001111000000111111110100001111010001110000001101110011110011000111011111111101111111111100010000010101000011110100001111000101110111000001110000110101000011001101010100110001000111010001001100110100110000111100001111000100010001000101111100010000000100010101110101011111000001110011110000000000000001110011000100011111010001110101111100,512'b11010101110100000000011101000100000011010101110000000001001111001100110101001101000111010001111101010111110011110101110101001101001100110111000011010011110111010101010000010000001100010000010111000000010000000111110101111100000011110100011111110000000000010101010011110000000001110100000000110101110001001100111100110100000100011111011100111100001100001111010100001100000001000100011101110100110111110000000011111111110001111111110100010000111100010011001101001111110011000000010000000101010101001101011100000000,512'b11001100010000001101010011001101110001010000111111000100001101010001000000000000110100010000011101010011010011000101111101001111011111111101011111111101110111110001001111110101110000000001110100010101000111011111000111111111111100000100111111010001110000110000111100000011010101001101000101001101011100010000111111110001110000010111000001010100000100000000000000110011110111000011001100011100110011000100110000111100010011000001000100011101010000000100010000000001011100111100110000001100011111001100001100000001,512'b01110111110100010000000101001100000011011100001111000111010111001100011101011101110001110001010011010111000011010000010100010101010011001100010011000000000101011101010001000111001111001111000001010011110000000100000011011111000000010000010101110000010100111100001100001101011101010111110111010101001101010001110000111100000111111101110011110001011111110000111111011111000011000000110111110000110011001100001100000000010100000111110100010111110000110011110001110101010011001101000100010000001111000000110011001100,512'b00010000000100011111000001010000000111010000000111010100000111000100010011111100000001111100000001000111000111000011000001010001001100010001000101110100000000011111001100010011010000111101001100111100110001110011000011001101010011010011110100001100000111110011011101000111000101010111010001000000110011000001000111011100010111000100010111110100110101110000110100110001001100110101010011110100110001011101000101010101000001110000000111000111110000011101110000010011110111011100010000111100001100110011010100000000,512'b01110001001101010000111111000101110111010111000101110001000011010000000101000111010100111100111111010000010000010101010111110101001101110000110000000001110000110111001101010000000001001111001101010100010101000100110011010100010000000000000101110011000111110000110000010000111111111101001101010100110000110001110011111100000001000111110011110100001111000111111101000111001100000101110001000000110101111100010111110001001111111111011101011111000001010111000111000001111101000101010001000100010001000011110001010100,512'b00110100010011010001000111001111011100010001001101110001010000001100000011110100110111001100000100000100010100000100000001111101110000110011110000010011000100111100111111010001011100010011111101110000110011010111110001000100110000000101110000111100010000000000010000110101010100010000000111000011110001001100000011001101001101000101000011000100110111011101001101010100001100010111001101000001000001011101111100011111111101110101111111000111000000010111000000000000111101010000111101110001010000010100011111011101,512'b00111100000011110101110000001100010001110100000011111101000111110111010101001111110100001101000100110100000101010101000011001111000111110100010000000000011100001101111101110000000100110011110111111100111101001100000111000000011101010100110000110111011100110000110000000111011111111111010100110111110111000000110100010100000001000101000101011111010000010101010011111111010001001111001100011100000100001100000100000101110000110111010011110011110101000100000101111100000011110000001111010011001100010011010100011111,512'b11111100000111111100010111001100010100110101001111000000000001010101110111000001000000010100011101110111111100000011001111000001000011010001110011010100000100011100001101010100010111011100010001000001000011110101110001000000000101000111010001000011000100111100001100111101010001010001001111001100110000111101011101110000111111000000110011110100110100000000011101010011010100111100011101110011000111001101011100111111000111001101111100110001010001010000000011010011110001110000011101010101010100000000000111011101,512'b01110001000000000011111100001100010100010101111100110001000011000011111111000011110000110000001100011101010001010100000000010100010100110100110000110011001111010111010001011101011111000000010000001111111101010001000011000100000101000101010011000111001100001111011101001100010000000001010100010100010000011101000100001101000011001101010001000101000000011111000101110111000000010001000101010011010100111111000101011100000011010101110111011100110101111101001100011100110011111101111101001111000011000101011100011111,512'b00001101000011110011110001000100011111010100010011110111000011110000000101000001001101110000000001001101011100000000010001000000110001110000000011110001010101010000111100010111110001000100110000010001000001010100000000000011110011010100010011011101110001000111000111001101000011111111000100000100111100000000000001000111000011110111000111001101000001000000000000110000110000110111010111010000000000000000110001111100110001010001000111111101010101010001010011111111010101110000000100010111000100001111010001110100,512'b11110000000001000001010100000001001111110000010001010001000011000101110011011100110011001100000111011101110011011101110111000001111100000101110111111101010111000100111111111100000000000001001101000000011100001100000000001100111100011101011100011101010000111100011101001111000000010001000111010101000001000100010011111100000000110011000000000000011100000000110111010001001111000001000001000001110000010001111111001101000000110011000001010111000011000001000001010100110000111111011100000111111101000000110011111111,512'b01111101011101111111011111010111010001001111011100110001001100001111000001001111000100010101010100001101110101011101011100111101001100010001011100000101001111110100111111011111000001001100001101010000011111000011110000000001010000000100011101000101000011110100010111010100010000001111011101010001000000010111000000110001000011110000000101001101010001111100010000000011000100000001110011110101001100000101110001010000111100001100000000110011110100000000001111010011000111011111110000011101110000110101111111000001,512'b11000111000101010001000011110000011100011101010101110101000011000000010001000000111100011101010101001101001111010000110011111101010001110001110000111111001101110111001101010011000001000001001111010111111101010000111101110111111100011100110101111100010011000100110001010111000011001100110011000000001111000000000001011111001100010100000100001111000100110001111111001111001100001100111100010100000011000101111101000011000001111100011100111111111111010111111111010000000101000100110100111101110011001100000100111101,512'b00010001000011011111000000110001011101000111010111110000000100010011000000111111000001011100000000110111000000000011010000110111110000110101010000110000001100000000001100011100011101000111011101000011000100011101000011010011000000110011010100110000000111010100010100000000110101001100110000001101000100111111000111000101010101011101000111010000011101000111110100000000110101111100010000000000111100010000010011000001110001010101001111010111011101110000000000010011110111010111110101000101000111010100111100011100,512'b01010000010001001100011111010101010001000111110111001100001101011111001111110011001111000101110101110111110100000000000001000011000011000000010011001111010001000111000000000000111111010000010001010001011101010011111100011101000001000001001100110001010000111100011101010100000000111111000011110111110111110111111100000011110111110001110111111100111100011101111100001101110101110000011100000100000011011100110100110101110001000111000100010101011100111111010101110001000011011101010000010011010000010011000001011101,512'b00110000010101001100111100111100110011110011011101011101010001000000000001001111110000000001000001001100000011010101000100000111010100000000000111011111000111110111001100110100001101011111010000001111110001111111010101010100010101000001000101110011010001000000110101111100010011000011110001110001011111010001110011011111000101000000000000000011010000010000110001011101010111110100110011110001110000110011110000001100010100010001000101000100001100010100000100000000010001011101110111010001001100011100001111110100,512'b01010101000001010100110000011101000001111111000011010000010011010011011101010100111111010000110101011100110100011101011100111111010001000111000111010000010100110101000001110011010100110101010000010001000101001111110100110011010111000101001111110011001100000000000101000100001101000101111101110001110000011100010101110111110011000000000101110100111100001101010000110001110000110100010100000011011111010100110100000001110100011111000101000111110111001100011101010001010001110000000000010100110101110100000000110001,512'b11110011010000001111000000011101111100011100000100010100000000000100110101000011010100110100010100111101000011000100010101011101000100011100001101110100000100010101011100001101000000011101011111110011010000001111011101111100001101110111001111110001110101000100000001000011010011000000010011000011000000000000010100011101000100011111110001000100110111000001011101010001010000110111110111111111000011111100110000110111110001110100001100110000111100010111110011110000011111110100000011111101110111001101000000000000,512'b01000101010100010000010111000000110111000001110000000111010101000100110111011111000101010011110001001111010001001100010000110101111111010000000100000001110100000100000000010101001101110100010100001100010000001100110001010111000001111100110001110000001100010101011111010011010111010101010000110101000001000111000000001111000001110101111111010000110111111101111100010000000101000100110000000101010101110000000011010100000000010001110101010011010001000001010001111101001101001101000100001101001100110001010001111100,512'b11010011110100110000011101111100010001111101111100110111011101010011111101110111010001010001111111000100010001000001000000000000010011001111010100000011111101011101001101010011000100011101000001011100000100000000000011000000110100010011010011001100001101111100000100110111010111110111110000000100001101110011011100000011001111110011111111111111110111010100110101011101001100010000000000010101110001000101110111000000011101011100000101110000000000110000111111010111000100000011011111001101000000000000111100011111,512'b01000011110101000011110111000011000101001100110000000011010100010001000000111101010011011100111100000000000001010000010011000111000100010100110001010111000001001100010001011100000100000111111101000000001100000101110111000111110100110001110011110001000001010100110000000011000100000000110100001101010000001111111111000111010000111100111100000001010101011100011100000000011101001111001100011111010011110000000000111111000000001111010000010111010011010000000000001101000000000111010100110001010101000011000001010000,512'b11110011000011001100010111110011111101001101010100011111010001000001000111001111010111110011010100011100110011110000010111000001110001011111011101110101000000000011110011000001011111010000010001000000110001111111010000110100010101000100111100000011110011110000010001110000010100000000000000000011010000111101001101000100010100111101010101110100000000001100111111010001010100011111010000000101000011000000000101110000000101001101000111111111110101010011010101000000111111000111010111010100010001000011110001111100,512'b00010101110100011101011100010101010001010001010100000001000000000000001111110100110000011101010001110101011101001100011101110011001111000101010111010111000100010001110000000001110011000011000100110011011101001111000101110101010011011111000000000111011111000000010000110001011111000011000000000111001111110001010001010000010000010111110001000001110111111100001100110111001101000101001101000101000101001100010100111100110000000011010100010101000101010001011100010101110000000111000011110000111100000011000100110011,512'b01001111010111010011110000011100010100000000111111000111000100000100000011000111000000011100011100110011110000011111110011010100011111111111010000000100000100000011000011000011000001111101011101010111010101000000110111001100010100011101011100110000110000001101010100010101000001010011000101000000001111000100110111000100111111000011111111001101110001010000111100110001011111010011110000110011000011010011011101011100111101010001111111010000001111110000111111001101010101000000000011000101111111011111010001110011,512'b00000101111111000100000001110100000001111100110011010101000000010000000001111100011101000000000011010000011101010000010101110000000000001111000001001100000100000011010011001100001101110111001100001100110100111111111101111111010011110100011101110001011111001100000000001111010111110100000100111101010001110011010011110101111101000101000000110101011100001101110001001100001100111111110000000100001111000100110000001101011101011100000000110000010100001111011100011100000001000111110100001100000101010000110101110100,512'b00110111010000001111000000111111110000001111110000001100110000011100110000110011010000010101000011000101000011010111000001000101110000011100001100001100001101011111001111110101010000010001110111011101000100011111010011000100110100110000000000011101000100011111110011010000000111010011010000000001010101111100111100001100110001010111000011001101000101010001011100110011011100111101010001110000010111010101000000010001111100111111001100110100011111001100000001110011010011000101000100110111110011111111001101000000,512'b01010111110001000000001101111101110000010011010111011100010001011111000101000001001100000100000001000011000011000101001100000101110100011111010001000101000000001100000000001111000101000000010111111111010000110011010100001100001100010001000000010000110101110111001101010101010100000011111100001100010011011100001111111101000111110001001101011101110100110101110000001100000100001101110000000000011100111101110001010100110101000000110101110111000100110101000011011100111101001111110101010101000000110100010000010001,512'b00000100000001011111000101000000011101000100010000011111011101010001010101000011011111110000001111110000111101000000010101110001010111000101111100010011000111110001110100011100010101000111110111110001000100011111010001000100110011010100110100010011011101110001110001010111010101000101000111110000111100110100000101110101010101110011011101000111110000110100010101000111111100011100010011000100000100111101111100110000110011001101011101010101010001010000000001111111110011110000011100111100010000001100111111010000,512'b01011111110011110101001101110000110101000001110000110101010100010001000011111101111100010011000111000000111111011111011111000011110100000001001100000100111111110001000011110001110000000111000100000111110100001111111101000111110001011101010001000101010100110111001100110101111101000111010011000011001100111111001101110000000000000001000001000000111101010101001111000111000001010111110000010111010000000101111111000101000111010101011101110000000101011100110100110000000101001101001101010000010011010000010111110000,512'b00011111000100001101010001010011000100010111110101010101011100110000000000000100110100111101111100110000110011010111110100110111010011000111001101000011110011001111111100010011010011000000111111001101010101001101011100011100000111000011110100001100110101001101000100011111111100000100000111000001010011010001000101011111110001000011111101110100111101110100000101000001010100011100011100110111001100000011010001110000000111010111011111010011010000000100001101001101010000001111001100000100000101110000010101010100,512'b00011100110000000000010100110000010001001111110011110000001111001100000101000011001101001111010000111111110101110001000001001111010011111101010111011101001101110101000011010011110011000100110001001101000011010011110011111100000100010011001101110000111101010011011101000101110011010111001100110100000011000101010111111100111101001111001101010101110000010011110011000001000101000111000011111111000011110011010100011111111100001100000001111100010001000111010101110101110100011100110011010000110000001100010001110011,512'b00111100010101111111010101000000001111111101000100001101000011001111111100000001000011110100110011010011000000111101001100010001110001000101110100000011010011010101111101000000110101111111110100010001000100001111000100000100001100110001010111111100000011000001111111000111010011010011110011110000110100000101011101011111000000110101001100001100110100111100000011010000110111010100110001111100000000010011010100110001000001111111110111110011000111001100011111001111011101001101110001011111110011000111000011001101,512'b11000000001100111101000001110000000000110011000011010111111111000001010101110001010111110000010101001100000000000100110100110101000100000001001100011101000100110111010111000100010011110011000100010001110000110011011111000011000011000000110011010100000111110011000001110001111111111101000011111100000101111111000101111111010011110011111100110001010000001101010101000101001111010111000001010000001111000101011101011111000000110001110100110000001111011111010011001100011101110111010111010100001100001111010001011101,512'b01110100010001000111111101000011011101110000000000000100010100000000001100000111010011000100111100111111011111000101000011011100001111110100000000011101110111110000111100000101110011110001010001110101001101001100011101110001011111000000000101000011000000111100110101011111110000011111011111000000001101001100001101011100110101001111110100000111000111110100010000110011010100111101000100000100010001000001110101010100000100000101111101000111001100000011110011001111011111011100001101010001110000011100111100110001,512'b11010000010100010111000111000001110111001100000000001100010000000011000100000001110111010111110111000000110001000100110000011101011111001101001100011111110011111100001100000101010100110101001100011100010111010100001101010000010000110100111100010111111111001101000111001100011101010101001100000000001111110000000001010100010011001100111111110100011100111101001101011111110100011101010101000000011111110101010111111100000011000001110111011100110111111101000000111100110001010101000011010000110111110011011101000000,512'b00000011110001010001011101000100010111111101000101001111110111001101110100011100000001000000010000010100010111110100011100010001011111111111111100011100011100011101000101000001011111110011000100000111000001110101110100110000110011110011010101011111000011110111000011011101010101000100000000110011011101010100110111001111110001110101111101001101000111111100011100001100000111010100000000000001000000000000000101110111000101110000110101010100000000000001010100010111000100000000000000111111000111000101010011111101,512'b00111111110000111100110101111100010011111101111100010101110111010001000011010101001101011100110100000100010001000101001100010001010000111111010001010001010100000001111100111100011101001111001100110000011101000101010000010011110101000101010111110101010101010011000011000101001100110100000000010011001100011100110111000000110101110111010111001101111101000000110111000100000000001101111100110100000011011111111101001100010101110100110001000000011111011100001100111111110011001100000101001101001111110011001111110111,512'b00010101000011000001010101011100011100110100000000010100110111011100001111110001110000010001110011111111110001000001011101111111000000010100111101010111001101110000110101001100000000110101111111110100010101110101000000010000110001011111000100110000001100011100111100000001000101010000110100001100010001110101011111011101110000010101111101111100111101011111110000111101011101111100010001011100110111010100110011010001001101000101000001000101000111111111011111010011110011110000000001011101010001000111001101000100,512'b11110101010001001100001100010100000001010100010001111111111111000011110100010000110001000100000011001111011111110011010100000101011101000111110001000100001100010001110011111101000000010111010001110011010011110001010100001100110111110100110100010111011100000000110011010101010100011100010000010000110011010100111101110000110011001101001100001100010101000001010011110011000100000000010011110100110001000001001111010101010100011101111100010011010001010000001111110101011101010011111100110000000000001100111100000111,512'b11000011000100000001011100000000000001010111010000011100111100110000011100010011000101000001110100010000110000000111010101010011111100110100110011110000010101000000000101000000111100000101010011010101110101000000010000010100010100010011111111001100110100010101010000000111000101110001111100010000000001110011110000011111000111010100110101010000110011000100000000110111110111010000000011001100010111110101010001010000010100110101010001110100000001010101110001000011010111010100110011001101001111010000011101000111,512'b00000101010101000001001100110100001111000100000000001111111100000000110001001101110101110011000001010011110000010111000100110111000001010100010001000011010111000000110111000101010011001100011101000111110000000101110011111101111111000111010100000111001100000111000011010000000100001100010001110000000000000111001100110000000111110100001111010000010001110000010011001101110100111111010011000001000101001111001101010000000001110100010111111101110000000001110000110001000101000000000111110101000101010000110011000000,512'b00011101000100001100110111000001001101011100000111010000000101001111000111010111000011111111010100000011001101111111110011010011010000010101001100010101000001010001011100010011000111010111000011000000010001111101011100000011110101010001111100110111011111011101000101111111000100000001001111000011000111010001001101111111000100000101010101010000000111011100000100110100010000001111000001010001000100110111110001010001010111001101000001011101111111000111010000001111001100110101110000010001010000010001111101111101,512'b01110011010000001111010101001100010100110100110111010101000111000000000011111100011101111111010000000100010011001100000011111101110111010100111100010101000000010101011101110101111111010001110111010101110000001100010000011101000001110000001100001101010000010111111111000111110000000000000000000001000000000011000111110101000100000001010100000011000011110111010011010001000011000011001111000111011101010101111101110000000011110001001101000100000100010100011101001111010111011111010111000001010000110111000111010111,512'b11000001111101001100000000110101110001010000000101000100000001010000111100111100010111110001110101001111010000110000111101111111001101110000000000000100001100010001001111001101000101010000110100110101000011001100110101011111010011000001110111000000010000011100001111010001001100010100001101110001010100111101110001000000011111010001110100000001111111000011000100000011010100000101010001000101000011110100001111110000111101110000010001011111011101000001010011010101110001000100111100010100010000000001000011000101,512'b00000000000101010001110000000001110001011111000100001111110001110101001100110001011100001111110100111111001100001101111100000101110000111100001101110011000100001100010100110100110111000101010101010111001111000000000000111100110001000100111101010000000111010111010101010000110011111100110100001100110100000100000001011101111111010011000000111111110011010111010111110101000111111111010000000011111100010111010111001101000011000101110001010111000111010000000101001100111111000000001101111111110011111101010100110101,512'b00110000010001000101001101111100001101010100110011011111111100010111000100000100111100000101011101000000010100011111001101111101010000001101010001000100000001000000010001000011011111011100011100001100010000000011110000110000010001110001111101000001000000001111110100000001110101010011011101111100110101110001010000001101000101011100010111110001000100000101010000110100111111010000000000110011010001010011011101011101000011001100110000000101010011110001111100110100010001110011110000001100000011010001010100110001,512'b11010001011100001111001100000101011111010001000011011101000111110001000000010000001100110011011100010000000000000000000100000011010001110101010111010011110101011100110011110001110111110111110101011100001100000101010101110001010011110111011101010001010111010001001101001111011100110100000100011101010101110000010111010100001100010111000001010011000100001101010011000000001100010100010001001111000011011100010101000001110100011100010011000011001100011111010001001101110011010111111101010000000011000011010000001111,512'b00000100000000000011001101010111000100000100000011000100110111110011011100000011000011001101111101001100010100001101001100001100110011000000110011010100000011110101110111011101000000110111001111000011011100000000000101000100110101000100110111010000011111010001001101010001001100001100010111001101110001110001010001110100000011000000001101110011110101010000001101111100011111110001110000010101000111000000110101110111011100001111010001010000010011000011000000110111110101110011110100000100010011111111110000010001,512'b01011111010111110111000001110100010101000101110011000000011100110011001101000101110001110000001111001100010000010000010011110001110011010101010100111111010101000101000000000100000011000011001101010001000000010100110100010000011111010100110011000000000100010001010100110000010000111101111101011100000111000101000101011111111100110100000101000011000011000111111100000011110011000100001101000011010100010000110111010000000000001111010101010011111111000001010011000001001101001100011101011100110011110001110001110001,512'b01110100111111010100110101001111010000011101000111010011110111010000010111011101110000000000110000010011110101110001001111110011111101111101110100110100011111111100110100001111010001111111011111001111010001111111011101000101010000010100000001000011110001000001000011000101110101111100000001001101011101000011000001011100110001010000111101010111011111010111011100010001001100011101010001011101011111011101000111000111000111000001111111110100111100111111110000111100010000001100001111011111000011110111001111111111,512'b01110001001100000111000100010000001101011111111101000101010000110111110000001111011100001101001111001101000001000100110101000011010000111101010100110000001101110001011111110111001100001100111111000100110000010101010111010000010100010011010000010011000111001100110001001111010011011101001100000111110111111101010011010101000011110011110011000101000100110000000101010111110000000101000000110001001101110111010011010011000000110001110101011100010111110111011111000111000000010100110111010101010100111111010001001111,512'b11010011000100000101011111110011110100110101010001010001000011010101110101010001000011010100110000000100111101010100011100010000110101000000110000110111000000111111111111110100000111111100110000010100110100000100010001001111110001010011000100011101000011011111110111000111001101011111011100001100110111111101001100000001000100010001110011111101001100011101000101000000010101001101001101000000110011011100011101010011011111000000000100010101000111000011111100010101010100010101111101110101000100110011111111011100,512'b00110011110111111101000011000000010001111101001100010011110000010111001111000001001100000101010001111111110000110000111100011111010001010001111100110100111101000001110001010100110011110111110011000100001101110011000100110001011100010011000000000101111111000000010000000100000011111101110000011100000011000000110101010011010001010000110100011101110111110101000011000100010011110101000000001101000011110111110000000001110100010000110011110100111100010000110000000000110011010001011100000101001111010001110101010000,512'b00011101110101111101001100010111010111110001010100001100110100010100110001010011110111000111001100000000010111011111000101000100110101001100110000010001001100111111110001110100000100011101111100001101110000000100110100110100110111011111010001000100011101110001000100000001000001001101001111110011001111001100011101110100110011000100111111010100000100001111110101110011111111000011000111000000010100001100111111000011011100000100010011000000110000011111000001001100110011110011110011011100010111111111000001000011,512'b01111111110000110000111111011111010101000001000000010100110000110100000111011101110111011111000001000100000011001100010100111111000111110000110011010001111101111100111101011101010000011111111100010111110011110011010101011100010100011100001100000001010001110000000001000000001111010001010011110111000111000100110000111101000001010101110111110011010000000011110111111100010011000000110001000011110011001100010000010000011111011100000011110000010101011100001101110111010101110011000101010000110111110011010000000100,512'b11001100000101010011000000111111110100001111110100000111010011010001010111110100010000111101110101010001110011000011111111001111011101110100011111000001110000001111010101110011011101110100000001010011111111111100110001000011001100011111111101000101001100010001010100010101000001010001110001010100001111110101001111110101000111000111010101110111000100000100010001010000110011010101111100000100111101011101010001000100000100011100010001010000000111110001111100000011110011110100011111110111010101000100010000010100,512'b01110101000001010100000100110101001100010011000100000000010001111111010111011101001101011100110001000001010011111100000111011111110100010100001100011100010000111101010000111101111100110011000111111101110001010001110100011100110011110011000011111101111100000011001101000000111111000011010000010011000000110111110100011111000000110100000011011100111100011101000100000011010001010111110000001101011100001100111100011100110001111101001111010101010000000101111101110001011100011111001111010111001100110100010111110001,512'b00011111010001000100000000110011110011001101010100000000010011001100011100010000010011010011010000110000000100110101110011011100001111111111011100110101000000000011000000000100010100001101111100010100111111011111000100111100011100000100110001001111001100010011110000000101001100000000011111000001000011001100001100000001000000010011110100111101011111000101010111000011011111000101001100000100010001010100000100000000001101110100001101011100000101000001000101000101000001111100111101010011000001001101001111110101,512'b01000101001100010101011100110111010111011101000111001111001111000000110001010000010001110001110101010111110000000001010100000101001111001111001111000100111111000101010100001111011111110000110101011111110111000011000100111111000100010100001101000111010100000100010100010000110000000011000100001101001101001111000100010111010111000001011100010001000011110111010100111100000000000000110011110101001111001100000000000100010100011111011111110101010101110100111111001111000100000000110011000100111111001100001101010011,512'b00110000000111010111001111000000110111010100111100010100010000000100010000110011011111000011000111010011010111010001010101010000110011110011000011110111110001000011111100111101011111001101110100000011010011000001000111110000000001010001110000110100001100110100110001001101001111011100000100011101011100010111110011000100001111110011110111010001110011000100010100010011000111011111001100110000000000110000110001010001000011011100000100110100010101000001110101010100000100010001000101010011000001001100110000001101,512'b00010001111111001111001101110101000111001111010100001101000100110011000100110001110101010011011100110001000001010101011111011101110001000111000101010011110001000111110001000001010011000000010011110000000101110100110011010100010111110011001100010101001111010111110101011100010101010001010001010000001100111111011111000100001111110111110111011111011100001100001100001111000000000111000101010011000001111101000011000101000001111101001100001101111111010000010001001100110101111100011111111111111100000100010100110100,512'b00110100110000010001110101111100010100110100010000110100111111111101011101010011000011010101010000011101010011001100010001010000000111110011110111010001111100111111000000001101111100000011110001001111010100110000110111000011001101000101010000110001010100000000000001010100000000001100111100111101110100000101011111110000010011110111010001000000010111111101000100001101000100111111010011110001001111000101000001111100011101000111110111110001010101001101110000000011001111001101011101010101010101000011111101010001,512'b00010100111100000101010111000101011111011101010011110011011100011111110001000111110011001101110100000001111100110011000011001101111111000001000001001111110011010111011100000011010001010100010000111100000000111101110111110100001111010011110011001100010111000100110100011111001111110111000011110101000001000011011100111111010100110001110111111100010111111111111111001100000111000100111101111101110000110100000111110111010000000101000001010000110101011100110111110000000000010100110101110101110100110011011100001100,512'b11011111010001000111110001110001000000010101010000000011110111110011110011001100000100111101010011001101000100110001110111000000000011010100001111110000010011000100111101001100010101111100001100110001000111110111111100111101000011000111011100110011000011110100010001000101011100001100110001001111111111110101110100110101010111010011000111010100010000110000110001000101000100110100011101110000000101110000010001000101000001111111010100010001000001000000110011111101000111110111010000001111000001001101001111110101,512'b11110011110001000111000101010011010111010011000100000100010100010100000000010111001101111100011100110000110011001111010111010111110011000001001100000001110011010101110101000001001111010011000000110100010000110101011101000011111111010101010000110011010100000101000011001100110000000001110000001100000000000111011111000101000111000101000011000011010011010111001101000111010011000100010011111100000000110100110101111100000100011101111100000111000000000101110000011101000001011111011101111111000100000000111100010000,512'b00110000000100110000110011000101110101000001000100011101010001000000110000000000000100011100111101001101001111111111110011001101000000000001010100001100000000010101010111000111010100010001011100010000001101000000110100000100000100111111000111001100000011010101000111110100010101110100001101111101010101010100110000000100010111011100110000010001110011001101010111110000110101001100111111110011000111000111110011001100110101010011011100110001011100111101010100000000010111000001010011110000000001110000110000110111,512'b11010011000011110001010011000111110011010111000001111101000011001101000001001100011100010001000001000011000111110011010001010100011101110100110111000011111100110100110100010111110001010111011101110011000100000001000000010000000100010101011101111100000001110101110111000001111100011111010100011101000001011111001111001101000100000001111111000111000000110011011101001101000011011101110111010100011100000000110001110101001101111100000100111100010111000000001101001101110001111101111111000100001100000111000111001111,512'b01000011010001000111110100110101110000111100110100111100001111000111110000000001110101010111001101010000011100110001000100111101010011110000011101000000110001010000001100010001011111110000001100010000010001000000011101110011110001001101001111000000010111110100010101110100111101000100000101001101010001110000010000011100010101111101001101111101111101111100111101000111010001001100111100000101110000011101000100000000000011010001000000111100001111000000111100011111000111000111010001110011000001111111111101000000,512'b00010101011101110101000111110000010000001101000000110101000000110100010011110111001111010001000000111100000001111100111100001111001100000100000111001101111101010100010000000101000100110111000100111101000011000001000111000101001101110100110011010100000100111100001101110011110100110100000111000011000011000000111100000001000111000000010011110111000100110101010111001100000100000100011100000001000001110111011101000111011100111100110011000001010101001101011111000011011101001101000000110001001100011100010000010111,512'b01111101000011111111011101000001010011000111000100011100110100000011010111110100000001011101000001110111001101110100110101010111010011000000001111001101000011010011011111111100001101001101011101110000001111111100111101010001110001010011111101111101110101111100011111001100010111011100011101010001011111011101000000000011000100110001010100000001010000010000110011000111010111000011010100110100010100011100000011110111110001001100011111011101000100000011000000010000010000001101110011000000010001010011001100000111,512'b01000100011101011101000100000001000100000011011100001111001100011111111111111111000001000101010101111100110100001100111100001101010101011100110111011100000011010101010100010101000011011100110111000111010000001101011100010001000000111101110000111100000001110101000101110100000011001111110011110001001111010011001100000111000111110111011111110001110001010101110011110100010011010001000100011101000000111101000001110000011100001111011111000000110100011111110100010000010101000101000111000011001111000100000000110111,512'b00001100011111010000000011010100010011000011000011011100001101010001011101111100010100110100000001110100010011001100000100110001000001000101010100011111011101110011000001011100011100011111011101010101000000000000000011000101111100011111110001000001111101111101010111010001000111000100110001111101111100110100000001000101010000000101110011110000000001000000010001110011000100110101000111010101011101110000000011110111010000110101111100010000010011111101110101000101001100010100001101000100110111000111111111000111,512'b00010000110100000001000001010111001101110011010100010100000000010011110011010000111111011100000011010100010100001101010001010100010100110100010111000111001100010100000111000011010001001101110101000100011100110100111101001100111111111101111101000011110011010011011101110111001101001101110000010000010011110100111101000000000001011101011100010000111111110000111100000111111100000000000101000100001100001100011111000111110100000000010001000100111101010000110011000101000001110001000100000000011111000011110100110001,512'b00010000001101000100011101111100110011010001001100000101010001000101011111010011110101000100011111110011000101011101010100000100000000000111111101000011000101110101000101111100011111111100000000011111000000010000000000000100011101000000110101011111000000000101000111111100000011011101010011010100010000010111111101011111011111110000010001000000110111011100110111000000010001011111011101010001010101010111010111001100000000110001110111011100011111010001111111110000010100000100001111010111010100001111111100010100,512'b11010100011111010000011111000111000001010101000011000001000101001101010100110001111111111100111101011101010011011100110001010000010101111100001100010101010011000100111100000101111111000001000111001101110111110011010000111101010001010000001101010100010000110000001101010001000011111100011111000011000100000000010000001101000111110000010000111111000100000001010000011100011101001111111100000000110100000011000000010011001101000100000111110100001101001111000100110111111100110100001111000011111111111111001111000001,512'b00001100000000001111000100001100110000110001110000111100000000110100111100000001010101000000001111110000000000000001010100011100110111110000000000110111110100110101000001001100110100000000111101010101001100111100011101010111001100000001001100010000110111000011010001110100110011000001000101110001110000001111110000111101111101110111110011000011000000000000000000010011000000111101011100001111000101011101111100110111001111001100001101110001001101011111011100110001001100110100000001000111111111011101011101000100,512'b00011100010000011101110101001101111111010111011111000100010100000111000001000001000000110011001101110100110000010111110000111101110000000111110011110000001101111100010100001100110011110101010100111100010000111100010101010011000011111100000111001101110100001101011101010101001100110011010001010001000001000001111111000111111111000000001111001101111100011100010001001101010111011111010001000011000100000011110111000000011100010100111111010001010101000000010011000000001100000000111111011100000001001100110011000111,512'b11000101010000111111010100010011000000000001000101000101000111110000110001110000001100010011000100110011110111011101111111000011001100010100010011110101110101110111111100001100000101000011110111001111110001110100110011110100010111110000000001000101010001001100001100000000010101000000010100111111110000010011000100000100000111110000000100010111010001000001011101000011000001011101001101000111011111110000111100011100000011110111000011000101001101111101000111001101011111010111011100011111111111010111111111111101,512'b01110111001111011111110100010000000000111100001101010100001100110100000001111101000111010011001101010011010011000001000001111100000100000111010000000000011101000001110011010000001111010100010111010101001100001101010001010101000000011101010001011100010000111100000100010101001100010000000011001100110100010011111100000101111101000100110100001100111111000100010000000000010101000001111100110011010101001101010100000101110111111100010000111101000101010101000100110101110011111100001100000000111100000000110011000101,512'b11010000110101001111000101111101111111001100001100010011111111000000110111110001000000110111011101000000000100010001011111010011001101000000000111000100001111110000000001111111111100010100010100000001010001010100001111001100110101010011000000000100011101000111010101000111110000000000010000000000000100010111001111111100110100000011110000111100000011001100001100011111010001011101000100000000110100000000010100010001010000000001001101111101000001010100010111000000011111010111111101110000110101110101010001001111,512'b01001111000001110000000100000000111100000101110000000100111111001111011111000100011101010011000011001101001100010101000000010100011101000100011111010001001101110100000101111100001100010111110001111101010000010011001111000100110000111100000111011100111101000011110100000011110000000000011101000100110100000000010011111111011100110100110001000101000001000011010001010001111101010000110011000101001100001100001111000000000100010000010101110000110000001101110100000101110011000011000111000101111101000000010011011100,512'b01010011000101110000000111001100000011011111001100011100001100111100110000011100110001000011011101001100011111010011110011011111010001110111001100011100011101001101001101010000000011111111010100000001110000000111001101000011110011110000111111001111011100001111000101000100001101110000000000010001110001000100000000111101001100001100011101000001010011110001000100010101011101010111000001011100010101111111010100111111001111001111010000011111110100110100000100110111011100001111110001001100010001000011000011010000,512'b01010001000101001111000000000001010001110100000100000000000100011111110000110001111111000001010111000000010100000011111100010000000000001101000111000011011101110101010111010001001101111100111100000100110101110011010001111101001111010100111111010100000111110101000011010111001100010001000000010001111100110111110001001101001100110101000001110001011101110101001111110000000011000100010100110001000111110100010000010001001101000000110111001100110111010000010000111100000001001100010000110011001101011101011101000001,512'b00110100010100110001000101110011010111110011011100010111010101010101110011001100011111000111010111000011001111111100010011000111110000010000110101000101011111110100010000011111000001010100000000000000110101000111000011111111000100001100000001011100010111000011110101011100000000011100110001000001110100010011110100001100010000001111000001011111000001110011110000000000000011001111000111110001111100011101000000000011110011110001111100000111110011110111010100010000110101110011110011001101000101110011111101001100,512'b00010001001111111101000011000101000001000101001100110111010101010100110000110011011111110111010001000011000000011100000111010011110001000011110111000111011100001100111100110011000000111111001100001111000011000000110100110100001111001111011101010100000101011100110000111100011100011100010001111100010111000100001100000000010111011101111101110111000001110100000000110000000111000011111111111101110100010000000000000100000111110101011100000111011101111111010000001111000100000101110101000000001101110100110111110100,512'b01000101001101110100001111000001001100011100000000110000000000010000011100011111000001110011010011110000000111010100001100010000110100000101010000000001110111001101001100000011111101001111000111010100010100011100000001001111110000001111110111010111000001010001110011001111010100110100001100011111111100010111000011001101011111111101111111010001010101010101001100010011010100011111011101010111000011000101001101110001110001110011000000000000111100011100110000110001000001000011110100000000000100000000010011010001,512'b01000100010011000000010100111100010001000100000101110011001101111101111111010100010101010100010001011100010100000101011100111111010100000000010111010001110001011101110000000101010101000001011100010101111100001101111111001100110000000101010000000111011111010000000111011111000100010111110111110100000000110001111101111101010000111111010100010000010111001101010101000101110111011101010101010111010111110011010101000001011100110011010011000111010000110000000001111111010100010000110000010101010101010000010011010111,512'b00000000000000110101110001011100001111010000111100000101000000110000110001010000010111010111110000110011010101001100111111000101011111000011000000110011000101010000000000010011000100010000000101010100110000011100010111000011010011010001110001001100000011011100001100001100110101011101010000010001000000000000010101010000000000011101001100001100010111110111011101000001010000000101110101000100010111000011001111000100110101110011010000010000000001001100110111000001110000000001111111000100010001001101110001000111,512'b11111100000000010101010101010001000000010100001111111100000101111111000101010000010011000111110100000001010000000001110101011100010011011100011111001111110000110000011111000101000001010100110001010101111100010000110100010101010011011101000000110111000000011101000111000111010101110011110100011100110001000101001101111111011111010000111100111100000111010011110001011100010001000000110111011111011101010001000111010011010011000011000011010101010000000111110111010101000001010111111111010000110000010011010011000000,512'b01110101001101010001011101000000001101010011110001000001001101111100111100000000000101111111000001000000110011001100000011111100010000000000011101000100011101000000111111001100010101010111111111010011110111110111000001110101110101000111000100000111110011111111010111000101001100110011000011110001110101110011011100011100000100110000000101110001001100110101001101000101000011000111010000010001001101110100010100111111000100110101010101000011111111111101000000000011000100001111000001110011110001111111000100110111,512'b11010111000000110001110101001100010000010111000001010100000111010100010011000100000011000111000011010100000011010100111100110001111100111111010100110001110101000111110011110000010111000101001100110000010100010111010111010100000001111111010000010100010001001100111111010101010100011100000100010111001111110011111100000111000011000111000000110000111100010101110001110001001101011101010000110001110000110000000100000011000100000011111111111100011100010101111100111111011111010000111111010101010001110000010000000011,512'b01110011110100000000110011000001011100011100000101111100110111011111001100110101010011000100010000110011110001110001110011000100110111000100000101000111110011110011010101010101000011110000001111111111111100011101010001111111110100010000110101010001011101010001000000000000010111011111010101000100000001001101010100111100000101110101010101010000110101010111001100000011110100000101110000010000110000011101111101110000000000000011000000010000110001111100111111010100000000010001010011110000001100011100010100001100,512'b00110111000001110001000111010101000101011100110001110111001101111111010011000101111101001100011111010000111101010000111100011100110101010001010111000101010111000100000101110001000001000111110001010011111111010011110100000000010100000011111100011100011100001100001101110001010111110101010111110111110001110100000100001111111100011111110001011111000100010101010001110100111111000111010001001100000001000101000100001100111100000011000011000000001101011100110011000100010000110100110001011100110101001111011100110011,512'b01000100010000110100010000010001111111110001001100001100000101010111010100010100000101111100001100010000111111000100110011001111110011010011010101110000001100010001001101110111110101000000010111001111000000110011110000110000000000000000001100000000001101010001110101000000000000001101011101011101000011111111111111110101001100000000110001010100001111010000000100011111000000000111010011010111010000110011000101111100110111000001110011000101000001010011010000000100000000000011011101110000110011000111111101110111,512'b00001101000011111111010111001100000011010001000101111111111111000011000001110001010011110011000100000000001101011101010100000000000001111100110100110001110100111111110001000111110001000001000000010101000101010100001101010011110100110001011101001100000011000100111101010101010011000101110111011100011111010101110100110111110000110000111100111100010011110011000101010011001100110000110000111111000101010000010001111101001111000101001101000100001101010000000111110001000100110000111100110001011101001111000011010111,512'b11111100000001110000110000010101111101110001000101000011110000000011110111110101010000000111010100010101010011000011110000110000110001001111110011000000000001010100000000010101010000110000001100000000111101010111000000000000000100111101000011010011011100010111000001011100011101000100110011000101110000001111001101010011000101010000000011110011110000110111010111110001000011000111010100111101110001000000000011110101000000001111000000011100010000010011010101110111011100000001000111001111000011110000011111010011,512'b11010011010100010000111111110011110011011111111100110011001111110100010101011111110001010100011111110000010111000111110001010011001111000011001111001101110111000111000100010000010101010101010011011111001100000100010111111111000000011100001111000000110000010011001100000000010100000100000000110100000001011101011111001111010111010111000111110000010100001100011111000001011101000011110001001100111111111100011100000000001111010011111100111101000001111100010111111111110000001100011111000000110011110000011111001111,512'b00000001000011010111010001110101110000110011111100010101110101010101000101000001010000000000000100000100011101010000010100010011000101011100110001001100010101010101010000000011000101000000000101001111010101110101110111000101110111000101110001110101010001000111001111010111010101111111110011010011000111010000010000111101111111110100010000110000010000111100011101010011001111001100000000001101000111000101000101111111001100010011011101010101110000110111010000010011110101000000000001011101110000000001000100011100,512'b01000011010000000011000001010001010000110011000111000100010000111111110000010011001101110001000100111111011101110100000001000011010101110000010111010001011100010101000000000001010000000000000100000001000001010001110011011100000000001100010100000000000111001100010011000000000101000001011101011100111101000000110001110100000011111100111111011101011100110111111111110011010111110100110000010000110111000101111111010011000011110000010100110011000011011111000100011101000111010111111100010100010000010100010001010100,512'b00000001110001010101110011111101010100010011110001110001110111111101110100111101011111010001001101010101111111110100011101011111111111111100110011111101000100000000110011010101011100000100010001011100111111110011001101010011010000110101000011011111010000110101001100110000111101110101000001010001011100010101010111010111110101010000010011110000111100000111011111001101010101110001001101011101110001110011001100110100011101110100000101010001111100000101000000110111000111011100000011001111011101000101000001110000,512'b00110001001101111101110001010101010100000100110011011100001100111111000101110111110101110100111101000001011111111101000101010001000101000001001101000100010011000101110111011101111111001100001100010000111111000101111101000101001100010100111100110011111100110001000100011111110101010001000000110100110101010100010001000000001111110000010001011111011100010001011111110100111111110001110100000011010000010001001101001101111111110011110001000101000111001101000100011111010011001111011111110011011101000100110100000111,512'b01011100000111000111011100011100000111010100000001000100111100011101110100010001000111110000010000010001000101110101000101111101010000110000000100111100000111010100000000000100110011011111001111010011011100010101110001001100010011000001010000110011001100000101110111001100110001110001000001000000000111110100000000001100001100111111010001111111000000000000010011010001010100000000110100000100111111000001001100111101000011010101001100011111001100000001110111110100111111000000110111011111110000000001110001010111,512'b01000011111101010011111101000000111100001111000101110111110101011100110011111101010101110111111111110001000111001100001111110000000000010000000100000000010011110001011100001111011100010111110011111100111100001101111100110111010100001101110101011101111100110111111101001111110001110100011100110000000011110101011101110100001101110111000100110100000100001101010011001111110111110100111111110100000000010000110001000101011100000011000000110101011100010011110000000111000000010100110000010000001100110111110000110001,512'b11011101110001110001001100000111000000000100110011110101010011000000000000110011000000110001111101000001110000000011111101000101010011000100001111010001010100000101010011011111110101001101000111110001010011010011001111000011110100011111001111010011110000110000010111010100001101011111001101110011010101110101110011000101110011111111110101000011000001001111110100000000110000000001010111111100000001000011001100000001010000010100000101110000000101000001110100011111001100000111000101000011010011110011000100000111,512'b11000011010101001111010001110000001101110001110111010001010101111101000011110100000100010100000100111101000100000000000100111101000000000011011101000001010011000001000101011101001111010001011101110100011100111100110000000111110000000000000011000000111101111101011100111111000011000011111101110101011101000101001111001111110111001111110011011100010100010000001100000111110000001101110000110011011111010011001100010101110100010000111101110100011101111111010101110011010011001100010101110000001101110000110000000111,512'b00000011110111110101000011000000000101010001111100010011110001001100000000001101110000000101010100011100010001011100000001010011000111111101110000000000010100110001000111000111010001110001010001110001111101000100011100010111010100000011011111110000010111010000010001000101011101111100010100010100110111000011000111000011010100110001000000000101010011001111110100010000010101000101010011001111000100010011000000011100010101110011011111011111010011001100001100001100000100110101110111110100011101111100110000110011,512'b00010001010000110011011111011111010111110101110100010000110011000100011101000000011100110000110111111101111111110100110100000011000001010000011111110111010111010011111100110101010100011111111111110111010100010101011111010111001101011111010111011100011100001100000011000001011101110111000000010111111101011100111101000001000101110001001111010111010100110100010101000001000011110001000001000100111101001101000100110101000001110001000011000111000011110000000100001100110000111111110001010100011100000100000101000111,512'b00010100001111110001001100010001011100011100011101010001010011010000110000011101000000000100010001010111011100000011111111000100010000110000111101000001000101000101110100010100000101111111010100000000111100011100010000110000010100110011110111000011001100110111001101110011000011000101000001000011000001001111111111000100010100010001010100000001010000000111001100010000011111010111110101111100001101110011110001000111110111000000010000110101011111011100110000010100000001110111011111000111010101110011011100011100,512'b11000111110100000011110111000011010111010000000001000011000000011100001111000000000000111111010000110100000101010011001111001100000111001100010011010100010111001100111111110000001101000011000001110000010000111100010111010101000111110111010011000001011101000111110000000101001100110111010101000011111101110100010100010001011100110101110011000111000111000111110100001100000100000111010111000000010011010101010000010101010011000101000000000001111101000111011101110101000111000001000011000100111100000101000111001111,512'b01000000000111000000110111110011110000010000110111001101001101000100110111110000110000000001011111011101001100010000111111000101110011110100010000110101000101010000110001010000001101001100011111001101000000111111111100111100110001010101001100110011110100000011000100011101110100010100000000010111110100010000000101000011011100110000001100010111110000110111000011010001110101010100000111110011000101011111010100110000010000011100010011000111010000011101111100000011011111000100110000000100111100000001010000000011,512'b11011100110101001100111100111101010100010100001111011111111101000001001100111111111111010001010100010011010101011111010101000100010011010101110101011101110001011101000000111101111111110011110001001111110100110000110001010111111101000111001111000011110000111100110000000011000000010111010100011100000001010101000100000000010001011101011111111101110000000100010100010100110101000111011100000000000101000100110100111100110001111101010011010101001100110111000011000011000001010001010101010011000000111111010001000101,512'b00011101111101001100000000010001001111000001010001000011110111010111111100111111001100111101010100010001000100110101010101000000000101010101001100000101000100110100000111111111000001110001110100010000000101000111111111000011110000110000011101010000110101000001011111010101010101000100110111001100001101011101001101110100010011110000110100111111110100010100010001110001110111110000001100110011010111010011111111111100000000110111111111011100011100010001110000000100000011010000010101000100011111110000110000011111,512'b11110100111100111101001111000001010101001101000011001111001101000111000111011101001111111100000001000011010000011111010000000100110100010101000100000000001100000111110111110101001100110111010100111100110101000111011100010101001111000011110111010111010100010011011111111100000111000100000011001100111111111100010101111101110000000111000011011101000000111111001111000000110101010011111111110011111100001100001100000100111111000111110011001111110100000001010000000011010001011101000101001101010000011101110001110001,512'b00000101111101000000000100000100011111000000110000000111000111001111011111010011001100010000000001010111110001111100010011000001011101000000000111111100000100111101011111010100001101110101000100000000111111000000011111111100110100011101010111110101001111000000001111011101000000011111000011011101001111000000011101000100111111111111001101010101000000010101110001111101010001011111010100110101001111000101001100010100000011010001110001001111010001110000010011010101111101000000001111001101000011111101010001000100,512'b11010011000000111101000111110000001101001101000001001101010100011100111100000000000000000000110000110011001100000111010001110000010100111111001100110001000001011111110000000001000111011100110111001101010001001100111111111101110111000000001111000011010001011100011100110101000101011111011100000000011101000011000100111100001111010111111111111100111101001100011101001111000111110000001101011101110111000000110100001101000000000001000000011101011111110000010101010011110101000101010001001111001100001111010001010011,512'b01010000010000010000001101010001010100000100000111000111110000110011001111010001010000010111010100011101110000010000111100000100111111000001110101001111010101000011000101011111010100000001000100110111010000010101011111000011010100000011001101010111010111011111110001010001000111001100010111011111000000000001000100001100110000110100000001000100000101001100000000000001010111011111111100001101001100010111010100000111110000110000000011110001011100110111011101011100001101111101000101111101000001010011000100001101,512'b11011100111111011111000000010001000100010001000001010111110011000000000001010101000011011111011100110001111111000000010001000000001101111111111101110100110100110100000011000001111101000100010100110001000000001100000111010101110111010011001100000111000101011111010000110011110011110101000101000111110101000001010001010011110000001111000111000001000100110011000100000001001101000100000001010000010000110000010011010001000001000111000001000100110011011101011100010111000100010100010000010101111100010000000101010101,512'b00110101000101000000010001011111001111110000001100110111001111000100000011000001110100111101000100110001000100000111010011110000010000001101010000001100111100110111110000010000000011010001000100110111011101000111010101010000110011001111001100110001010001111100010001000001110011010101010000111111010101000100010111110111000011010001110000000100011100001101110011000000001100000101110001011100001111011111010001110000010001010011001101110011000011110001010100010001000111000000000001011101001101110000110000000000,512'b01111100001100011100111100000111001101111111110000001111010001011111000001010101000101110001110011011101111111110011011111111100001101000000110100110000010000001101001101110000110101000111000000110000110100001101000101011100010101111100001101111111011100110011000000010101011101001100000101000000010001001111010000000011001100110101011111111101010100000001110100001101110001000011110000000001110001110000010100000011011100000101110111111101110101110111001111000101110111001111001100010111110000110111011100010101,512'b11110101110001010000011111000001110100010001000100010001000001111111110100001100011100000000110111010000001101010000001100000000110001110111001100000001110101001101110111111111001100000011111111110100011111001111000000000000110101110111110000000100000000010111110001010011110000000101010011000101011100000101001111111100011101110001000011000000010000010100000000000101000011000100000011001100000000001100001100000000010111000100000011000001110011110101111100000001110000110101110000000100000101001101010111110100,512'b00000011110101010111011111001111010000000111001101111101000100000101000111111111010101110001110100000011111111001100001100111111001101010001110000010000000111010100010000110001111111010111000111111111011111010000110100001111011101000001110000000111001101000100000001110001110000000111000001111111000100110000110011011100011101010100000000001111010011010111000001001101010101110111001100001111000011010101010101011101000001010001110111001100011100010100000101111111001111000001110100010111110100110001000001011111,512'b00010011010111000111010100000011111111001100010100000011010000010101001101000001010001000001001111111100110111001100111111110101000001010011000011011101000111110100001100011101011101010000000001010111000000110000111100000000001101000001001100010000000101000100110000110000110111011101000000011100000000000111000011110011110000001111000000000001000101000000110000001101001101010111011101110000010101000011000101110100110111000000111111000001011111110001110000000011000101000101000101001101001111110111010111110101,512'b11000011000001110011010000110001010001011101110011000011111100010111000111010111110000010100110101000111111111010001000100011101011100110101000011110011000100000001010001010011110000010000010000010001000001010001001100001100110100000000010000111101001101110000001111000111010000010001000111000000000000110111001101000000110001110000011100110001011100110011001100010100011101000100010011010111010000000111011100010001001111000011010001110101110100010100111100000100110100010000011100010100000001110000110011010100,512'b11110100011101110101000100000000011101010011001100000111011111010000010001010101000000010100111100000100110100010111001101000011010100000000011100000001010101010000010101000101111111011100010011111100110001111100110000001100111111000101000011000000001100010001000100000011111100000001010011000000001100110000110111010100000011000101000100010000110111000000001111110100010011110011000111110000000011110001110101000011011111110011010011110100010100110111110001110101000100001101010001010000010000110111000000000100,512'b11110011011111010011110111001111110101000011011101000000001101000011000011010100000111111100000001001100110011011100000011110011010001000111011111110100010000010100011101010011010011110000110111000101110000110000001111000101111101010000110101110101010111001111111100111100110011000000000011000100110001111100001111001100010100000000110101000111001101000101001100000101001100110001000000110101000000000111000001000001000011110000111111010100000001011111000011111100001111000001010000000111010000111111110100110101,512'b00000111000001000101001101010101000111111100111111000100110101010101010111110001000111001101010111000000010001000000110000001101000111111101110111110000010101011100010101110001010011010001001101110111011100000000010111010000011101010011010001001100110100011101011111001101000011000111000001110100110111011111110100110101110100000011110101011100000000011100111100010011000011110000000001000111111101000101111100010000000001010011000111010000011111010111000101011100010100000000000100111101010000010101011101110001,512'b01000101010000001100010001010000001101110100011100000011000000110101001100110001010001001101110111111100001111010101010100001111010001010111111111111101110101010011011101110111010000000111110001111100111101010011011100010111011101110101010000110000000001110101010111000000001101010000001111001101011111001100000100010111111101111100001101110001000100000011001100110000110101111100110100011101011101011111110011010000110001010111000111111100011111110001000011000011110100110101000111110000000111111111000000000111,512'b01001100010001000100110011000101010000110001000101000100110100110101111111000011110011000100110000000111110000111101010001001100011111011101001111011111110011110100110011111100011100010011010001010001110000010101110100010101111101110101011111000001010101010111000011001100000111010000010001000111111100010101011100000111110101011111000000110000111101011101001111000111110011111101110011000100110111010111111111110011010000010111000111110100000101000000110011001100001101011111010100000000001100010111000100000101,512'b11111100000111010011000001010101111100001100011101010100010000000000000111010001000011010101110011000011001111010101011101010001010000000101010011011100000001110111110011000011000001001100000100000111110011000001000001000111000000000111001100010100001100000100111101110000001100001100011101001111000000110111010001110001010001011101000011010111010001010111111100000011000011110000001100001111010000010001110111111111110000010011110000011111001111010000011111111101011100011111111101000001110011000101110111000111,512'b01111101010001001111000100110000010000011101010011000000011101110011001101110011110100010111000011001100010000010001110101110000110000000111000001001101010101110101000101000101011111010101000101010101001111001111000011001100110101110001111111000111001111000000000011000011110100000000001100000001010001110100111101000011111111001101110101011111011111010101110000110000011101010001000100111111001101000011010111000111110011110001110011110101000101000100011100000011110000011101010100110101111101110001011100001111,512'b00111100001111011111000011110001000000110000001111011101000101110001000100011101011111010000001111010100110001000001010101000000011111000001011100000011010101110111010111010001011101001101110111000100010001000000001101110100010111010111111111010111000000010101000000000100110101110100000001000000110001110111000011000100110100000100010001111100010000110001111100110000001111110001110100000011010101000001010000000100111111000111011111110000011111000101001111001111010111110100011100110011110111000100110000000011,512'b01001101110000000001110111011101000100011101111100110000000111110001010000010100000000110100011100111111110111000000111100110101010001000100011101010000110101111101110100001101000001001101110101110001000011011101000111110101001101001100000011001100001111110001011101001111010111010101111101001111000011001100010001010001000000000100110011010100110011000001110000010001111101110000110001110001110011001111000100111100001100111111000000011111011101000111110101010101110100001111110001001101011101010100011101110000,512'b00000001010100010100010001001101000111001100010100110011011111000001010001010101000000000001110001000001111100001100001100010011111100000001111101000001110011000100010000111111110100010011010111110101000011011111011101010100111101010000000001110000110100000011000100000001010000000001000100000111000011001101010001010001010001110101000011001111000101110100110000001100001111001111010001001101011111010011010011000100001100110011110111000101010000010000111111011100001111000111000100110100010100001101111111011101,512'b01000101010111001100110001010100010000001100010101110011000101010000110000111111000111111100011111110011010101010001011111110011010000111101111101000001001101110011000001010001110011111101010101110000011101000001010000010001110111001100000001001100010101001111010000010001011101001111010100110101000000001100000000000000010100000000110100000001011111110100111100000011001101011111010100001100110011110111000001000101110101000000010111010011000000000011010000110101011101110000000001010011111101010001011100001101,512'b01010100000011000000001101000000010001000101110111001111000001010000110100001101110011011101010000110000000100110111000001001100000000011100110000111100111101110111110000110100000011010001010101001100110001110100001100110101000100010001010111000011111111011100001100111100110101011100110100110011110000110000001101011100000000010100001101000011010111001100110111010000010011001100110000110100011111111111111100011100001101010000001101000111110000011100000000000011010001110001000101010111010101110011010111011100,512'b11000100011111011100001101010011000111110101001101111100010101110100110011010111000101010001011101011101110100001111010011010001111111110111001111010000110011001101001111110000010101000101110001000011010011111111110001111111001100111101110101000000000000000001010100010100010011010011010101001100011100110011111101110100001111000111111111110100110001010001110011010100110001011111000101110011000111010101010111110100110100000001110011011111000000111101001111110001000000110000000000010000010001000001110100000000,512'b00000011010001001111110000011100110001010111010001010101000011001100000001010001000011110011110101010011010000111101011101000100110100011101111101110011111100000100110000010100111101110100010101111111110000110100001100011101000100000111011101110000001100011100111100010111110000010000001100000001110101110000010100010101010011000101010101110100000000110000011101000100010011000100000000110101010011000101011100000101000111000111011100010001010011111101000101110000110111001101011111111111110000010001110011110011,512'b00010111110001111100110100110111001100111101110100111101000101000100011100010100011101010111000001000100000011010011000111011100011101110000001100010100010000111111000111000100110000001111011111000100011111110000000000000101010111000000110100110100001111000101010011000111011111000011000111110100010011010000000111001101010001111111110000010001001111010000001100011101000111010101110101001100010011110001010111000001001111001111010001010101110000000000010101010001001101010001011100001111000011111101000111000000,512'b11001100001100011101110111010101000011110011000011010111000101110001000011000000011111011101010100000000010100111100000000001111011100111111000100111101110011110100010100000011110001010111000101001111110001001101000000011101010000011100110001000111011101011101010001001100001111110000001111010101001100001100000000001100010000010011010000110101110001011101110011010101010101001101000001110100000111000011110011001111011111000011111101010011110011001101111111010001000101010011000101110101111101001100111111110100,512'b11000011000001000011010100011101111101111111000011000111110001010000011111010000110100010000010101110001010101010000011111000001111111010000010001110001110101110111110100110011011100010001011100110011110001000111011101110000000111010111000011000101000001010100000000010001000101110011011111010011000100010101010100010001011100001100110000110011110000001101001101010001111111011101000000000111111111001111001100000001000001001100110001110000110000000000010000000000110100000000010100010000001101001101001101001100,512'b00110001111100001100010101001100010111001101110001011100001111001100110100010111110100001111000100001101000011000101010001110011110100011101010001111100110000001100010100110101110100010000110101010101110100110101111101011101110000000101010011110101000111111101011111010001000101001111010001010111110101000001001100001111111100010101010101110011111100010111000111011100011111010100110100000001001100001101000001000100110111111111110000000111000000110101000000111111011100001111010011110000110111001101010000110111,512'b00110111010101001100110101000100010111000100011100000000111111111101000011110100000001000000000100111101000001000000010001000000010000011100000011011100000100000000110001001111010101110100010011010100110100011111010000110001010001000000000100010001001100110000110000010111000100111100000000011111110001011100001111110101011100011111000101010000111100110000111100011101010111110000011100011101010100110000111101110000011111011100110011000011001101111111110001000000011111111100000000000101000000010001111101001111,512'b11110000110111010100110101110111000101110000000101000111010100010111000101011101010101110101110011001100010011111111010000110000110101001101001101000101011111110011000101000101011100000011010100110000110000011111111100000000000000110101010000010111110000000111010000000100111100001100110000110011000101010101110011000011010111110001001111000000011100000011000101111111110011010101000001000011011100000101000000000101000001011100011111000000111111000011010001001100001101110111011101011101000000011111111101000100,512'b00111111001101011101011101111101000001110011000011110011000000011100010000111111010111001100010011011100001100010101110100000000110111110000010000010100010011010000110100000101111101010101110101110011110001000000011100110111110100010000000000010000010001001101010101110100110101010000010001110111111101000111010111000001110000011101000001011100000100000100010000110001001101011100001111000011000000110000000101111100000100110101000100110000000100010000110001011100000000111100001100010111000100010001001101110001,512'b11011111000011000000000001011111011101110000011100000100000011000100110100000000010100001101000101110101001100000001010001110111110001110001000100111101010011001111010111111101001101011100000100000100001100000011000011110001010101110001000101010111110101000011000011010011110011000101010000000000110001000100010111110011010000110111000100000000010001001111110011011101010011111100000001110100000101011111000011000011000000001100000001010100110011010100000011000111010000000100010100111100110001111111000000011111,512'b01000001011100000101000001000000010100010000000001010000110011111100000001011101010100110000110000010011000000110011011111011111110000011101001101111111010001001100011111110001000000000101110011010111011111010011010000110100011100001100001101010001000101111100010111000100001100000100011101000100111100000011001111000011000111011101000101011111000011010011001100110111010111001101010111011111110111000101001111000001001111001100010101010011000000110001001100001100010001010001000011000100010011000100110001010101,512'b00110001110000001101000000001100000100001111111101110011000011000000111100000000000001111101011100110111000011011100010101010011010101011100111100001111011101110100000100010100000100110000000101110000010011000101110011001111010001111101111100111111111100110101110000010011010001110101000101111111110111010000001100010001110101001111110100111101110100110001111111111111000101000101000100011111001101110011110100000100110011000100010101111111011111000100010001000100001100001111011111110011110101001100110100000001,512'b00000000110011001111011100011111010000110001110000011101000100110111010100110101010000111111010101111100110011011111010101110000000001000000001101001101010100010111000101111101110000010001010101011101110011000001001101000100000100010100000011110001111101110100001100011100111101000000110000010000010101111101010001110001111111110000001101000001010000110000000001000000010111010001010101111111010100010001010000000000110001000100110000010000001111110011010000110100111111000001001100001100000001111101010000111111,512'b11010000010001010101010111111100000000110000000100010111110100001101111101010100000100000000010011000111011100000001110100110000110100111101111100110001010011010111011100010000110101000101001100000001010000010000010100110000000000110011000011110100110011010001110011000000000100010001010011110011001101001100010111000111000100011101000101000111010100111100110011110001110011011111010000001101111101010111010111001100111101011100111101000001010100010100000011001100000100110111110011000011010001110011001111000101,512'b00001100000100110011010011001111110000010011111100000100110100000111110011110011001111010011110100000011111100001100011111010001110001110000010111001100011100001100010101111111001100010111110101111101010101110101010000000100111100111100011111000111111111000000111111010001110011110101010111000111010001010101010111000100110101110100111111000101000000001111111111000101110011000011111101010011110111000100000111010011010001000100001100010000010100001111110000000000011100010001111101010001010101010001110101010011,512'b00111100011101010000110001010101111100000100110000011101010001111100001100000111000001110101110101110000111100111111000011111101110011010001010100110101111111110001111101111101110100000011000111000111001111010001000011111100010000000011110001010000010100110111000100011111000101110001110001000011111100001111010100110000000001111101110001110000110001011100110001111100010001110000000101110111011101010101000000111111000101010000110001001100001111010101110111111101010101010100010101010000001100001111110100010101,512'b01000001000111011101010011010001010100010101000101011100010101000100010111011101110100010011010111110011010000000011010001001101011100000011001100000001111111000101111100000100000000010011110001000000000001001101000100000100110000001101110001110000111100000001000000001111111111000001111111010011000100000100010000010000000000111100000001000100001101111111110001110011011100001100010011111101010000001100000111010000001100010101010001000000110001110101000100110100010111000111110101010111010000010011011111000000,512'b11110000110011011111000011001101000011000000000001001111010101001101000011000001000000010000011100001111010000111111010011010101000100000101000101011111000011001100110000001111111100111101000100010100000000001101011101111100010000001101000011110011011111000001010001111100010011000000111111111100111111000101000111110000001101111100010100000101110001010000010011011100011101010000111111000100010111001101010100001100000101011100110011111101110111010011010011000101000100111101011101010000010001000011000000011101,512'b01001100110100110100000111000001010111000100000111011100111100000101110001010001000001110000001111000011110000000000110111000100001100110100000000000011010100111100010100110011010011110011000011010100001111000001111100000100110001010000010011000000010000110101110101110100011100000001000001000011110101001100011111010111001101011100011100110001000001000011011101010011110011110111000001110101000100000001000001011101010111001111111101001101000011010100001101000100110101000101001101010101000011010000110111110101,512'b11111100000101011101000101010100010100000111010011010001110100011100011100111101001111010000111101110011010000000011001101110011110101010100110111000111010111001100011111000100011100000000111111010000111101110011110011011111110011001111110001001101000111010101011101000101110011111101110100011101000011000111010100000111001100111111000011000100010000010000110000111100110100011100010111001111011101010111010111011101010001000100010111011101000001110000010000010111000000000100001100110000010101001111010101000000,512'b01001111110100000111111100010011010111010111000101001111010101010100001100001111110011110001001101010000011101011100000100111101010000010001000001001101001101000000010011000011011101011100010001001111110100000001010001001100110001010100000100110001011111010111000101000011011101001100000111000101000101000100000100000001000000000101000000010111111100010011111100010100111111000101010100010101011101000001001111010001110011110001110001010101010111000011000100111100110000110111011111000001110000011111001101110011,512'b01110000011101010111001111110011000011000111111100001100111111000000010011000011000001110100010001001100011111111100000001110001110011001101000111000011010011000001110001110100110100001101010000111100001100110101110111001111110011011101010111001111010000010000111111000001111100001100011111000101000111110011010111110000000101000000010011000001111100110011110000110100000111110011010000011100010011001100000011111100000111110001110001000000001100000000010111000011110101110111000100111111011100010001110100010100,512'b00010000000001000100000000110011000000111101110111001100001100110101111101010101110101010000011101010100010011111111000101000100010011010000000001110100110100010000010101000111001111000011000001011100111111011101110000010001111100001101011101010011110101111100111101000001010000110000001111111111000100110001110011010101000011010001000001010000010111001100010100000000010001110011000111000001010011001101000101010011010011011111000001001111001101010111000011001100111100000011111111110001110001001100011111000001,512'b11110101000000111100111100110011011101110001000101110101001100000100111100010111110000010101000001001111000000001100011101011101000100010011010000011111000100110100011101110000111100001111010011111101010001111101000000011101010000000011010100001111001100001100000101001111010101000100000100000100110011011100011100000011001100110100110101110111000011000001001101010100110100001100000011110000001100111100010001000000110100010001010000001111110001011111000101000011010011001100000011110011000100010111010011010101,512'b01011101110111001100010100110000000101001101010001110011000001000101110011010011010000110111110000010011111100110011111111000001010000000111010101010001000011001100010000000011001100010100111101001100001101000011010001000011010111111111000000010101111111001111010101000100000111110000000101110101001111000100011100000011111101001101000011010111000001000100000001111101110001000100110011000001110011011100000000001101110100010111000001001100000001011111110000110101110111000111000001110001001100111100010101010011,512'b01010001010000011100110111010000110000110001111100000001000011000100000100110100110100010000110001010011110100000100010000010000000111110100000011010000010101001111000100010000010011111101011101110000000000110001010000110100000000010101010011000001001100110011011101011111011100011111010111000100000000110100110000110011110011001101001111000101010101110101010011011100011101000011000101110111111100010101000111000100110101001111000000010000110101110000000011000000110000000111000000000100000011000100111111010101,512'b00110011111101000111000101000000000011111111110100010011000001000111001100010000110001110100000100010111000001000111011100110100010111110101010100000011010100001100010101000001000111111111000000111100000100001101110011110000010000111100110101000000001101001111010000000100011111001100000000011111000101110000010001010101000011001111000111010000000101000111010101110100110101110011000100111100110000010001110001110111110001110001111101010001010100011111000001000101010011010011000111111111111100010011001101001101,512'b01110101010011000001010001110111001111000101110000110100000100000100000000000111001100110100000101011100011111010100001101111111110011010101010000110000011100011100000101000000000111110111111101001101000000001111010011010001010111010011010000110101010011001100011101010100000001110111111100110101001100000100010111011101011111110001001111000100000100110001110011111100000101111101000100000001000111001101110001110100000100000011001111010001001101000111001100011100000101010011000000010100011100000000001111010111,512'b11000000010000011101011100000111111100110100110000010001001111000101111101001111000000001111010001110100110111111111010111011100110100001100001100001111000111001111010000110100000101011100110000110000110011110111110000010100000111001100011100000100010000001100111100010011110101000001010101000000011111001100111111000001010111000111110001011111010100001101111111001100011111010111110101110101001100000111010100010100011100010100110101110011110111011111111111010011000011010000000000010000000100000011010000000001,512'b00001111111101110011001101010111000001000011010001001100011111010101010001011100110001110011011100110100111111010001010100010100111111111111001111010101000001011100011100001100010100000111010100010101110000110111110101001101110011110101110011000001110011110000111100011100110011110101001100000001010100000000010011010101110000010011010100000011001111011111010100000101110100001101110101000001110111110100010000010000111111001100000011001100110001000001000011001100010100001100011100000011000100000100011100110011,512'b00000001011100011111011111000100000001110101111111110100110011000001110100010001011100010000011101111100000001001101000011010000000100110111110100010011010100110011001101010101111100001111001111010111000011110000000011010011000011010111000000010111011101010000000100000000111111000100000100000000000111000111010001111100111101110011000101001101110100000101000101000101000111010100010011000100110001010100010100110101110100110001110011010011111100000101111101000111011101001100010001000001010111110001111111011101,512'b01110101010000010011010000111100111100010001010001001101010000010000000001010011000111110001010000111101110111010011000111111100000111111101011111000011001111110000111111110111000000000100001111000000010001110011011111000101010101110000001101111101001100011100111100011100000100010011010100110011011111110001000000000000110000011100110000010101010100001100110100110000010001010011000001010100010000000011010111010101110001110001000101111100011100110000110101001100010111111101010101010101011101000100011111110101,512'b00000001011100110011000000110000111100110100010100000001000000000001111100010000010101000100001101111100000101000000000011010001110101110111110001000100011101001101000001000000111101001101011100010111010101010011010101110011011100000101000100111111010001010011001100011101000000010000010101010001000011010001001111001101110101001101011101010100110011001100111111011101110001110111001111111111000111110111110111001101111101000001110011110101000011110001001101000101010100110100110011000000111101001100111101111111,512'b00000100010100000101011111010000010100010000000001000100000111000011001101000000110000110001000101110000110100011111001111111111110000011100001100011111000001110001010001010001110011000001010000001100010100010011010001001100110111010011000001000101001100110111111100001100110011000101010000110111110000110000010011000011001100010111110011111101010111000100110001000100111101110011011111111101111100000011000100110100110011010001000001000000000000110000000001001111110001010011010000000101010000110000110101010011,512'b11010001001111000000010011111101111100001100110011000100010001000111001101000100000001010001001101001100110100000011000111011100010001001101010000000001000111111101111100000101010000111100111100010101110000001111000101111111001101000000110001001100010100111100110111000100010000110101111111011100010100010000000000110100110101001100001101011100011111111101000101110000110000110011010100010100001101010111000000000111010011010100010001010001001111010011000111011100000001111100000000011101000001110000000011001100,512'b01111100110001110101000011011100111100111111111111110000110000010101111111010011010111000100011101110101111101110100110100111101011100110001111101000011011100001111000101010100000011010001010111001100000001010000110111010001000100010111110101111101000100000000000100111100001101000111011100110011000000000101010111110000000101010001001111111101110111000111000001110001000000011111010001010100110000010001000001000001000000010100110001000100110101010100011101011111011111111101110100011101000011110111010001000000,512'b00000111110011001100001100010000110011011101001100110000110001110001011101010101010101011111110011000011010011110011110001110011000011011101000111000100110001000100000100000001001111001111111101011100001101000000110000001101001101110111000100010101011111000011001111010101111111001111111101000011010100001111110000000001110011010111000100001111010111001101010111110011000111011101000101111100110001011100011101111111110001001100011100010011110111111101011111001100001100001101010001111101000101000101110001010001,512'b00010011000011001111001100000111000011111101010111001100000000000100000000010100000000010100001101000100011111010001110000111100010101000100000100011111111100010111001100000011000111010000000000111100000011111100010101000001110111110000000001010100000000001100010011111101110101000000110100111100000100111101110000000001001101000011000011110000111111000001010011000101110001011100000101110000001101110011111100111101010111001100110100000011010100110101010100001111010000011111111101110111000011110111001111000001,512'b00110111110111110000011100000001110101010111001111010100001100000000010011110100110000010100001100110011010001000000011111110100111101110101111101010011001111111111000100111100000000011111010001000101000100010000001100010001011100000000110011110101110011000111111111001101001111001100000100010011000100000101110001011100111101001111111101000000000001000101010000010100010101011101111101110000111111110001110001001100111100011100110111000011110001011100110101111101000100000100000101110100110011110000111100110000,512'b00001100001101010000010001011101000100001101001100010100110000111101110111000101000011010000010100000011110111110100000101011100010000010100000100000101000000000101000011001111000000000100110001110000010111011100011100000101000100110001010000000011000111010101001111010000110001010001110000000100111111110111000111001101000100011111000100010111110001011101001101010100110100001100000000010100010000000001000000110111110011110001010111010001000011111100110100000001000011011101110000110101110000011111001100000000,512'b11000100001100001111000111001111001111011101000100000101110000001111111101000000000011000001000011110001011111110001001100000001001101010100111100110100001101010111110101010011001111011111110100001101000011000101000011001101010011000011000000110101010011000111110000001101011101000101000000001101010100000111000100000101111100110111011100001101011101010100111111000011111101110001110100110011110000111111000111000101001101110000111111110100010001000100110101000001011100110001010001010011000011110001110100110111,512'b11111111011111111101110111000000111100110101001101001101000011011111000001110100010111111101010000000011010000110101010111110100000101010100000000010111010100110111000001000011011101001111001101110101000000110000010000110011011111000001010100000100110011010000111100000000010011000100010111010100010011010011010001000011110001011101000000111101000100000000000011110000110000000111010101111111000011010000010011011100110111010101110111011101111111000011000101110001000111111111000100110100001101011100011101000001,512'b00111101110011010001010011110000001111111111010000000001001111111111010001110100110011000000000001011111010001010101111101000101010001010100000111001100001111110011001100110001000001011100111100000100000101000100110000110001010000110001000000010100110100000111000101110001010011010100000011110101000000010101000100110000010001110111111101110000110100010001011111111111000100010101010001001111010100010100010101010100110011111100000100110000011100001101110000010001110000001100110000010111000000110011110000110101,512'b11001111001100000011110100111100110111110000000011000000010000000001111100000100011100111111010101010001001100000001110111000100010011111100000100000111010001000011000011110100111111111111010011000000001101001101000101110100110100011100001111111101000000001101010011000100000100000101010100110001000001110111110000110011001100110001110000000011010001111111110101110100111100000000010101010111000101010011010100110100110001011101000100000011010011000100011100010011111111010001000111010011000111011111001111110101,512'b11110111110000110000001100001101001101011101110100000100000011000001001101111111110100000001110000000100000101001100110111000100011101110100111100000011110100000011010000010100110011010101000001000100010100001101001111110101010100010011110100110001001111000001011101110101011101110101111101000100010111000000110101011100000100000101010100000100000001010100010001111111000111111101000001010000001111000011110011000000001101000100010101010000010011000000010001000100001111001100010100001100000001011111011101111111,512'b00110111000101001100110101001101011100001101010011110100010000010100000100110111111101110101110011010001001101001111000011010001110111000000000000000100010001000101110111111100010111000100111101110000110001000101010100110111001101010100110011011111011111000111001101010001010000010100001100011100110000000001011100000001000011001111000001000001000100010101000001111100110111110001000001010001001100111111110100011111111101110000000111110111010100110001000100010100000011110000001100111101000011011100010111010001,512'b01001100000000001101001101000001000011110001010000010001000000000111010101110100000000011101010011010101001111000100010001111111011100001111010101111100111111000111110111010101011100111111000001110001000011000011000000000000110001010100000000001101111101010100111100001101111100010111111111110011010001110100010001010000000100000011000001000001001100111100010111010011010000110001110111110000110011111101110011110011001111110011010011000101000001111100011111010101000101000000010001110111110101001111001111110111,512'b11011100010011111101001111010001111111011101000001010011000001110000011100010001010011010100010111110011000001110000010100010000001100000000001101001101110111110100011101010011000111011111110001010111010101111111110100010111010001000011000011010011010011010001010001000101001100000101010111111101011101000011111101000111111101011100000001000000111100000011010011010101010101110001000000111100000101111100010101000101011101000111010111000001000000000011011100010011110000110000010001010100000100010101010011110111,512'b01110100000100110100011101111101000011000001110011110011010001110011000101000001110000110001011101111100010101000001000000111101110000000111010111010000110011000001111101000101011100111111000011110001111100010000000000010100110100110000010000001100011111000101000001010100010000011100011111010001010100111100010100010001111111010001110101000101000101010100000011111100110011010000110000010111011101010000010101000100000001000011010101111101110111000011001101110100000011110100011101110101001101010001010000110000,512'b01111111001111010101010000110001000100110011001101000101000001001111010000110000110111010011000000110011111100110001010011110100000100000101001100000111010001110000001100010100110001000000011100011111110011000100010000001111110000110100011100110101010011000011001101110100000100010011010100000101000000001101000000110011000011111100000101010101111111011101000100011101010011110001010011010000010000000001010111111100110111011100000100000100000100000000010111111100010000000000000111011100110000000101010001001100,512'b11111111000000000011111100011100111101110011111100001100111100000101000011010101000011001100010001110001010001010101110100010000001101011111110000010011111100010001000111010100010100000011110111000000110000001100000000110001111100001101000111000001110111010100011101010000000001110000110000010011010101001100110101001111110000010011000011000101000011001111000001110000001111001111010001110111110011011111000100001100011101010100110000000000010001010111010011011111001101011100010101110001000100111100011100111101,512'b01001100001101110000000011111100010001110101111111010011000011001111010101000100110101111100010100000001010001000011111101010001010111000101010111001101000111111101000011001111000001010011010101000001000100010100010101110101000111001101000011010101011100010101010000110111001100010111001100010001001101000000111101111111011101010011001101110001000100111111000001000001000011000011000000011111000100110000111100110101110000000111000011001111000100110000110000010011001111010001001111110100000000010001000000111100,512'b00000011011111001101111111111111010000111101000000000100000001001101111111110000000000111111000001000000110000000111111101110100000101001111011100010000010101111100000101000101011100110101010011011101010111000001110011000100010001001101110100000000000000000011110000110100010000010011000001110100010100110100000101010100001101011100111101110100110101110001000001011101000100111101011111001101010001011100010100011111001100000011110011001111000011110100000100011100000001110000000011110101011100000100001101010101,512'b00001111010000010000110111110101011100001111001111010100110100110000011111000001000101001100001100110100000001110000000000110000001111011101110000010111010101011111000111001111110100010101010000010100000001001100010100110011000000010111000000011111110111010100000111010001010000011100111101001101110001001100000111000001011111110001010101010011110111001101110100000001110011010111010000110100001101000111110111110000111100000001000011011100001101110011111100011111000111110111010000010011010100010011000000001100,512'b00010000110000110001010000111111000011011100010000110011011101110011010011010100110001110000110101000111000100000111000111010111000011110011010000010100111100001100000101010100011111001111001101110100001100010001001111110111000100000101110111111101110100010001110000001111000111110101000101001111010111110001010001001100010001001101010100011100010001001100000000010100110001001101010100110111000100110000110000111111000101001100001111010111111100110001111101011101011111010000010000110101011111110111010011010001,512'b01110001110111001100110001110001011100110111000001000100011101010001000111010011000000110001010111010111010011111111010111000000000000110011001100110100011100110011011100110001111100110001010100000011110011110000010101110000000001001101001101110000110000110111111101110101000100110000000000000000010011010100010000110101110101110011110001010001001111000001011101110011111111011101110100010100010111000111110100110111011100010011001100001111000101111101010001110011000000001111111111110101110100110101110001011101,512'b01010100011100010111110101110011011111110111000111010101010101111100000101011101110101000100001100110111000001000111000111001101010101010011010101011101111101000011000101011100010001011100110000110000001101010001000111000011010101010100010000010111011111110011010111010111110000011101001100000000011100001101000000001100000100110100110011000111001100000100010001010101000101010100110101001100111100010001001101010001110011000011110001111100001101110100011111010111011100110100010011110100000011110100000100000000,512'b00010011000001001101010001010000011100110001010001000001000011111101001111011111110100010011111111010101111100000100000111000000110100001100000100010001010111010101011100010001111101010101000101000001011100010111000111000100011100111101010001111100001111000000110100111100000001010011001100000001111111110011110001001111000100011111110100111100010100010000010000001100001100110111110101000100000101010101110111000000001101000100110001110011010100011101000000110100000000000000000111001111000000110001010101110000,512'b11000111110111010101110101010011110011000011011100110101001111010000001100001111110000010100000001010011010100110001110101000011001100000100011111001100000011000100011100010100110101010000000100110000010011000000111100110000010001001111110001000011010111010011010011000001111100110000000011111101010001010100000100000111000100001100001100011101010000010100010001110001011101000100000000110100000011010001001101110000111111000100110001001101000001000000010101011111001100110011000111001111010001000100110101001101,512'b00000100010011110011110000001100000000010111001101110111010001000100110011011101110111110001010001000111001101111100111101110000011100111101000011000000011101111111010000000111010011110000001100000111110101001101110011010011010100011111000000110000011101111101111100010000010100000001000001011111110000111100110000000101111111000101000001000101110100000100010000110111001101110111111111010001110111001100010100000100001101001100110011010000000001000011000101110001000111001100000100000100000111000001010001000000,512'b00000000000100111111010001001100010000001111010011110001000001110111010000000100011101010101110001110001000111000101110100010000010011010001010100001101000011001100110011000100000011000101010000010001001111110101111111001100110101010111011101110111001111000001110001011101110111010000000001010011000100010001010100110001000111010001000000001100000011111101110011010001000000011100000101010100010000110101010001000111110001000001010011011100000111110011000001000000111111000111000100111111110000110000010011000100,512'b00110111110111010011110000000111111111000100011101010100000011111101010111001100110011110100110100010000010011010111010000110001000000000000000000111111000000111111010011010101001111110111010000000001110111010000110101010011110101110011000100010001110001000001010111111101010001001100110000111101001100010111010001010101010111010001111100000100000011010100000101011111010001011111111101110000011101110000000100010101110100000100000101000101010100010100110100110111110011010001010111001111110111110011111111110101,512'b00010100010111001111010000000100111111110001110001011101110111001101110000000111000011110011111100110000110000010100111101111101010100110001111100001100001101011100000000011111011101110011011101010011001101001100111100000001000111110101000101000101010101000001000000010011111100011100001100010011000100001100110101001100111100110001000011010000010000110011110100000000111101010111110001000111111101111111001100010000000011110001011100010101110000001100110000110000011111000001110100111100010011110101000111000000,512'b01000100000101010101110001001100111101001101110000001111110111110001001100111101010011001100110011010101001100011101000101010111000000011100010011110101111101110011000000110011110001110101110000011101000001000100111111001100000100000100000001011100111101000100011100010000001100001111000001110011011101001101110101000000110000000011111111010000000101000100110000010100000111000001110000000111010011111101110000000000010000001111110000111111110100010100011100010001011100011111001111110101111101110011000000111111,512'b11001101110101000001110001001100001101000011010111001100110001011100000101110011000000001100000100001101000011111100111111000101110011000111010011000101010000010100110011111111000100000011110001110101001100111111011101110100110111010000010011000111010001111111010100010111000101110100110100010000000001010000001111111111010011000000010100111111110001010111010011000101000000110100010011110111010100010101111100110101000011110000110011010000010100110001001100010000001111010000111100000011000011010111000101010000,512'b01110000000001010111110001000000001100000000000000000001011111000100111111000101001100010001011111000100000100011111010101010001000011011111110001110001000011000000110100011111110111010111000111010111110011000001011111000111000000000111111100000011000000011111110011010001010011111101011100110111010100001100011100110001110000011100000001011101010011110011110001110011001111000011110011000100111100110101110111010101000000010011110000001101000011000100010100111111011100000100011100000011010000110100010011001111,512'b11110101010011000101110000011100010011001111000100111100110111000000111101110001110001010011010011000111111101110000010000111101010000110111111100111111111100111111000001110100110100011111111111001111010111110000000000000100010001000011000001110000000000000011010011010111000111000000011100000100010101011101010101000100000101111101010100000100000000110100010101110000110100110111111100110000010000011100000000011111110101000100010000000001010100010001001100110000110001111100010000000100111101000011010111110000,512'b01000100000000011111011111000100001101110111001111000001110000111100010000000000110100011101000011000000010000110000000000000111010000010100000100000111110001000001010011000101010111110111000100000101000000000100110001010100011101001101010011000100110101010111001100011101110001000000010101111111011101010100011101010101000000010000000001000011010101000001111100110101111111110101010100000111111101000100110011110101000001000101001101110111111100110101110101000100000001010000011101111111001101010001000101000011,512'b11110101110000000001000000010001001100010001001111001100010011010111001100111100010000110100010001001100110101000000001100111111010100110100000001001111110101010011011100000100110011000001000100010000001101000100110000011101110111111100000100000100000011011100010011110011111101110000000000011100010101011100011101110000000011111101010011001111010101110000011101110011111101011100010001000011000111010000110000010000111111110011111101011101000001000111011100000101010111010100011111001101010000110111011100110101,512'b11110000010000000001011101011100010100110011111111010111111111000011000000110101010100010011010111010011110011010001110111010100010111010000001100000011000000000111010001000000000001001101001100110111000011010100001100010101011111000101000000000011011111110000011100110001111101000011000000110001110001000111110100001100001100011111111111110001010011001100000000010000010001110001000111010111010011010011110100110001111100011100001111110001000011000001000000010001001100110101111100001101000000000101110101110100,512'b01110000001101011101110001001100001100110011010101111100010000110011110001000001011100010111000001110001001111001101111101110111000001001101111101000111000101010100010111110100000011010000000001010011110011000100011101000000110100000101001100011101010000111111110100000000000001001101000000000000111111000101010000000011010011001100110100010001010100011101000001110101000011111101000111000000001101000001111111010111010001001100000001110100110101001100000111110100110000110100110000011100110000110100110000111111,512'b01010111000001001111110000000001111100111100000101011101001111000111011101110011010111010100000100110011000111001100011100000001011101111111000100111100010011000100001101000101111101001100000000111111001111110100110011011101010100001100000011001111001100011100000000000001000001010111000001110100110011000101110001001101000011110001000011010101011101110101110001110000111111111111000011010011000100000111001111000000010111111111000011110000001101000000000100011111011100110100000100000000010001000111110001110000,512'b00011111010101110011110011010000001101110111110011010001000000110001001100001100000001110000011100011111010101110111010111111111001111111101111101110111010000001101000001001100111101011111001111111100110100010001110000001101111100000001110101000111110011110111110101000100000001111100000001010011110111010111010011010111001111111100110100111111111101010011110100010101010011000111010011011100111111000100110100000001110111010001110100000101010100010100001111000001001111011101110100111100000011110011110001001111,512'b01011111000001010011000011000011010011111101000100111100110001010011010000010001110000010000010011001100000101110100110000000100011100111111111100010111000111000000000001010101111111001100001101110101110011010111010111000101001101000101111111010011110001000000000001110001000011111101010111010001110101010011000100001111010011011101110100001100111101000101001100110100001111001100110100111101001100010011010100011111111111000000110100111101001100011100111101000111010011001100010101000000000101000001001101000001,512'b01011111000001110111110011001101011100111111111100001100110100000011010000000001010100010101011101011100000101011111010000111101110101001100001111010111011100001100010101010001000100010011000100010001010101001111110011001111010011000111110000011101011111110111000011011101000000001100111111010011010011110001010111000001000100000001111100010001000100110111010101000101110001001100000011110001011101010000001101000111000001001111000011010001111100110000110000010100110101110000000000110111110000000111110011010000,512'b01001101010101000101011101110000000111000001110001110100001111110111001101010011010001110000110100010100010100011100111101000100000001110011110111010011010000010101110100010000001100010011001111000011010000110111110111000000110111110101000011000000110011110100000011001111001101111101010001011100010011011100110000000000010001010011000101110101000101111111111111010111000000110101011100010000000001000011011100111101011111010011110100011111001101110111011100011111010000000001010001000111110100110001111111010000,512'b11001100000001111101110001111101011101000001001111110001001100011111000100111111011111010001111100000100001100000001000101011101000100111101011101000011110001110111110100111100011100000011110001000011001100000100010001110111001111001101110101000001010011011111001111000011000000110011010001110111110101000111000100011111010111110000010001110111110011001100000000011100010101111100001111000100110000011101000100110001111100110111010000000011111101010100001101010000011100010000000001010111010000000111001101111101,512'b01110000000011001111011101000101011100110011111100110001000101010001001100110011000011110000110100010000110011001100111100110100011100010100111101010001000001000111110101011111110000011100001101001111010111001100110011000100110000110011010001110000110001111101000011000101010011111111010001000111110001110100000001110111111100110011001111000100000011011111111100000000000100110111000011110000010111000011110000001100000100110011110011110111011100011100010100000000111100111111001111000001000000110101001100110111,512'b01110101110001011100010000110001111100011101010000000001010011110100001111000100000100000000000001000101001100111100000000010100001111001111000011110000111100000000010111110011010001110011011100000011110101111111110001111111110100010000111101010011010100110011000011000111110011111111000101001101011111000000111111111101000100000100111101010101110000000001001101000111001100000101000000001111000001000111000001000001110000010001001100011100110111010011110000010011110100000111000101011100111111010011000000001100,512'b11000000000001001100000000010000111101011111001100011100110001110001000000111100000011000111111111000001011100111111001111011101000001010001000101000000010001010000011101000100001100010000010000010111001111010101010011000000110001110000010100110001110001010111110011010101010101110011000001110111011101110100010111010001110000000100010100000000110001000100000001011100010111001101000101110000110001010000000001010111010100001101000101111111010111110111110001110001110000010100011100010000000100110100000101001101,512'b00010101000000000000110001011101111101011101000011110001010000110001000100011111000000111101001101001111000001011101011100001101000000001111000001000001110011110011001100000100000111000011000000110001000111000011000000001100000000000001110011001111000100010000000101001111001101110111010101000101111100110001010100010001010001110000001100001100010001110000001100001111000001011100110000011111010011110011011101110100010000110101000111000000011101111100011100000001010100000000110111011111010100110011000011110001,512'b11011101000001001101010011010000001100111111010111010101000100000100010011001111110001011100011101000101110100111100010111000011000011010111010101110101110101000111110011000000001101110101001100111101000011000100111100010111110101010000110111111101011100110000000011010000000100010101010100010011010111000100110001001101010001001100110111110011110101010100000111000000001100011100010100000001110000001101110011010111010000001111010100011111001101110111000111011100110011011101111100000000110101010100110001010011,512'b11001100111111110001110100111100010111110100111111000101110001000111110001010111010000000100000100000001110101011101010011010011001100000101000101010001110101110011000011000000000101000000011111011101000001000100000000011111011101010001110111110101000100011111110011000111000000010111010111111101111100111101000001000000110000000001111101001101110100110011111111000001000011110100010100010000111100010001111100110100110111000000001101010011000000001111001111001100011100111101011100000000000111001101001111000001,512'b00000101011100010101001100000011010000001100000000010011011101011101000111000101110101000101010000011111110001110100110101111111010100001101010101111111000100110100010000110101110000000000000001010111000000010000000101011100010101110011010000110100000011010000111111110011110000110100000011000001000111010100011101110000110001001100001100010001111100110011011100110101110000000100001100010001010001110000010111111100010001000100011100000011111111110000000101111111011100001101000000011100000101110011001100111111,512'b00110000010001110100000000010000000011011111110011010111010000010101010011000101110000010000110101111111010101010011001101111101001101000000001100001101110011010000010011000000110001110101111111010000000111000001010000111100001100001101010000000100011100001101011100000001000100110101000101010011000000010011110001000011011100011101000100001101001101011101110011011101001100011101010111010000010101011111000001111111110000010001000001010101110101001101110100110011001101010100110001001111000101010000110000110000,512'b00001100111100000001010100000100110101111101001111110101000100111111000001000001111111111101010100010001010111001111110001010000110101000101110101110011010100000001000001001100001101000111001101010111000111111100000111010000001100010001001101001101111111110000001101011101110101010101111100110101110001111111010011000100001111000101011100001111110001011100000001001100000011110001010100110000110000010001010101110101110011001100011111000000000011110000010101010000001101000000110100011100000000110101010001010100,512'b11000100110100001111110000001111000001010111111100000000110001000011000111010111010111111101001111110100001100110111110001010101110000000111001100010000000001011100110111000100010000000101111100010011010011110100000100111101000100000000010101110011000001111100111100001100000101110011110101111100010101011101001101110000000100110011001100110100111100001111110001111111010011110111111100000000010001110000000001001100000100011100010100000001000101010000110101110000011111000011110001000111111101001100010011111100,512'b00010001111111000011000001110001011101010001001100000011001101010011110101110000010100010100110000110000110100000101001100010100010111111101011101000001001100000000011100111101110001000111001101010011000101000000010100110101011101010111110100010001010001110001111111010100010011000000000111000000000000000011000111010101110101001111011101111100111100110111000111000000000001001101110011010100000000011111000001110000110001010011000101011100111100010000011101111111011100110100111101000000010001111100010101110111,512'b11000101000011010011001100110100000101001111010001011100001101011111110000001111111101110011011111000001110011110111110000110000010000000100000111010101110000110111110000110001010000010100000100011100000100010011001101001100001101001111011100000100011111110011001101110000011101001111011100000000010001000001111100110000000111111101111100000011111111001100111100110001010101000000001101110100110000110101111101001101111100110101000101000100110000001101001101001101000001110101000001111100010111000001000000001100,512'b11001111000111000000110100010100111111001111110000000100000100010000000011011100111101110000000111110111001101010111110011000000000001000101001101110100011100111101001111001100010101110011000111001100110101000111011111110000011100110000010011000000001101111101001100111111111111010100010000000000010000010111011101001101001100110111010000110011000111011111000111000000111101111100010011010000001100000000001111000100000111000001010100111100010000000100110111010000001100110011110000001111000111000111010111110001,512'b00010111000000011101111100110000011101000100010000111111001101001101011111011100000100001111010000001111110100000111001100010001000001001111001100010000000011110001000000111100110001010011010011001100000100010101010000010001010111001100000000010111001101010000000000001101000111110100110011001111001111110011000100111111000011010011001100000100000111000100001100000001110000001111000101111100010000000101110000110001110000011100110000000100110001010111111100011101110111110100000101110011000101111111001101001111,512'b01000100000101001111010101110000111100010101000000001100110011010111000001010001010000000111001111000101010100010001011111010001111100010000000101110100010111001101110001000011111100110111000111011111110000000111001100010001010100000100001111010000000100001111010101010011010101110001110100010100111100110000001101110100000000110101001100110000010111001111010100111100011111110111010001010101000100001100110101010000000011111101000111000000010101001111111101010011110011000100011111111100110000111111111101110011,512'b01011111000101001100110111000000001111010011110101010011010001110100010000110001110011000100110100001101110111001111000101011111011100110100010111001101010111011100110101001111010001000101010001010111011100110011011111011111010100010100111100010100010000010111010011000100010101000111000000011101010000000011010111010111111111000101011101011111000000111100000001000101000011010100111100010011110100010111000011110100000100110011111100001111110000110100000100000011110111000100110111110100000000011100010000000011,512'b00011111010000000011000000110100110011001111010100000100110011000100010011000100011100010101001111000111010111110001000100010000010011000001000011011111000001000111010111001100001100110011110101000001000101110001110011000000001111111101000101111100011101010001010001000101000101111101010100011111001111001111011101110100111101010111010000001101110111011100000001110111110100111111001111010000110111000100110000000000110111010001000101110000011101001100010000010000000100000001010100110001001101010001111100010011,512'b00111101111100001100010000111100000100001101111101110101010111000001010011001100110001010000010100000001000001000100000000111100111111000011001111110101001100110101011111111101010001010101000101111100001111010001010001000000000101110011110111000000011101010000000011001100000100110001010011000000110111001100000011011111000001010100011101010000000101010011001100000100011111110000110001000001010101110100110011001100000111010001111101111111000000001100001100110000001111000000110001111101111100000101011111111111,512'b00010001010000011100011111000000111111000000110101000000110111010000000000010100000000110100000000000000110100000100010001111101011111000001111111000001011111010000000000011101001111110011000111111101110101000101000011000101000011011101110000010001010100000000000001011101000001010001011101010011110001010111001101110111000001000100000000000000110100010101110001011111000011000100000001000101111100010100000001010001000000000111001111010000000000110100001101110100010001011100000011000011110001010011110011010011,512'b11011101000101000000000001001111000000001111000101110001110011010000010001111100110000001101001101110001110111001111110000011111000000000000001111001101011111010101010100110000110000000101001100110101110100110001011101000000010100000111000101011101010101110101010000110011010001000100110000010001110011110111110011110100111100000001110011110000111101000100110000110111000100010011110111001111000001110100000000001100011111000011010000010111000000111100010011111101111100110111110101111101000100110000000100000111,512'b11000011010011000101001101001100010011000000110011000000111111110011010000111111000001001111000100000001111100110001000000110100010011110011110000000101000111110000110011001111010101010100010011111100111111000101010000110111111101001100010000110000111100000111001100000001000000110001011101110011001100011111010100000011110011010011110011110011111100110011110000110111111111000101111101000101111100000001000100010001010011000001010100000000110101010000000101110101111101110001000111001100000100000111110101011100,512'b11111101000100000101111101001100010011001100010011010100000011001111000011110000010101000111011111010111011100000111001101110000110111111111001111010000010100000100000011001111110100000101000011001100010001000011011111000001000101110001110001010001010111010111000001110001001100001101000100110001010101010100001111110001010001000001010000010001010011000100000000110001001111000001000011000011111101001100110101000111010100001100000001001100010111000001010111000000110100000001000100010011001101000111011111111111,512'b11001101110111001100110001110101110100000101000100011100110101011111111100110101000011000111001101000000010011010000011101000001010001110001010001010001000101010000110100000101010101011111010100001111000111001100000100011100011100001100110100111100011111110011111101010001010000000000110101011111000000010111011111000011111100000100010101000101001101000100010101110101010101010111000011001111010111010100010011000001010001011100111101110000001111110011000011110000000000110000110100110001111100110000011111010100,512'b00011111000101000111110111000001110011110001110101110000001101110001010100001101011100010000011100011101000101111111001100010011010000000011110111011100000011111111111101000000001111000001010000001101000011110100000001110100000011011101111100011100000101010101110011000000010000000101001100011101111111110011001111011101000001110111110000111100111100110111000011110011011101000011110101011111000001001100011100000000010000010100111100110111001100110001111111001100110000011101001111110101010111111111111100110111,512'b00110100110101010001000000001111000111111100010111110001010100011111000001001100110100000001010111110011000001110100011111011101011111110111000100110001000000000000000011000000110000110111110101000111010111001100110000010100110111000001000100111111110000011101000100000000010011001101001111010000000000000100110100011100000011000111110111111101010001000001000001010100110101110011000011000100001101000101010111110001001101010111001100011101011101000000111100011111110001000111001111110011110100000100000011111101,512'b00000100010011000000010101110001000101110000110011000101010100011100010000111100001101010000000100010100001111110011110100011111001101111101010001000011110011000011110001111100111101010011000000010000110000000011001100010100000001010000110011010000010100001100000011000111111101110000111100010111011100111101000100110001011100000101011111110100000100110000110101000001110000010001000011111101110001000100010011011111000011000101111100010011010111000001111111110100110011011100010101000000011100110011011101110100,512'b11010101001101111101001100110000010011000000010101010101001100110100000101001111111100111111010101001100110100001100000000111101000100110100000111110011110100011111010111000001011111000101000111001100110001111111110100111100111111010111110001010111001111110000001100001100001111110100111100000011110000000111111111000011011111010011000101111111010001010000111111010000000101010101110011011111000111111111110000110100001100000101110100000000110001001111010000111100111101110000110000111100001100010000110000110001,512'b00010111110100000001001101110011110111110000000011000101001100011100001100010011000100000100001101000101111100001101010100111101000100010011000100000101110111000100110111000000010000010100111100110001010011110101110111111111000100000111000011011100110000000101001111000100010001000100110000111101010111000101110001110100000101000011010000011101110001010100011101010100110000000000110011001111110111010011001100110011111100010000000111010111000000010111000001010001010011111100001100010111011101010011000100111111,512'b11000100010101001101110111110000010000110100000101001100000111000011110011010111110011000011011101011100000001011101000000110100000101000101000000010100010000111100111100010111010000110101010100110101000101110000000001000100000011000111001101110011011111011100011111111101010001110001010111000001000000110000110100001100010100000011000101110111010000011100000001010011010011110011001101111111001100000111010000110100011101000011000100000111010100111100110111001101110101001100001111110101111101011111001100110111,512'b01011101000000111101110001011111010100001111001111110101011111010100000111110000000101010111001111001100110011010000001100000000010100011111000100000011011100011101111111011101111100001111010000001101110011000011010011000111001111111111000100111100001111000001010100001100010011010011010100010111000001000101110011011111110100000001010000000000000000011100110001000101011100000100110000010100000100110001110100010000010000000011110111010011011111010111110000010100110011000101111100111101110100011111010011001100,512'b01110101000000110001010100000111010001000011000011010000001101000011001101001101010011010000110101010100000100010011011100010100010100000001110000000001010001110100010011010011000101110000110001110100110100011111010000011100110100110011010011110001110001010000010100010011010011110111110011010011110001110011010101111100110000010001000000111111110100010000111100000001001111000101000100000100111100000100000001011100111100111101110101010000000000010001000100110100010000000011110011000001000011000111000000111101,512'b01011101011111010011011100001111110011001100111111110101110000001100010000000101110011000100110011011111010000000001000000000100000000000000000101010101111111000011000011110001110100000011110111110100010000111111011111001111000000011111110101111101000000010111110111011101000101001101000001111111010111000100001111010111000101010001010001010101010001000000110111000101110111110101000100111100000111000000011111001101011100000011001111001101110100011111000000010100000001001111110100110001001100111100000001000000,512'b01001101011101000111010100011101111101111101001111110100010000000101111100110101000101111101110111000011010101110011000100110101011100110000010101000100000111001101011101011111010100001100011111110011011100000111000100010000000001110000010000010011000011000000110000110011111100000101011111000001001111000101011111010001110100111111011100010100110111001111010000111100011101010001010000110100010111111111000000010000000111000000110100010000001101010101010111001101010011000100111100000001000101000001000001000000,512'b01110001000001000101110000001101010100001111010000001100000000110100000100000011001100011100110111001100001101000000010011111100000101000000110111111111010101110000010111011100000011010001110001010011111100110111000011110000001101010000110100001111010101001101010101011111111100110000000101110111001100011100110000010111010000110000000001010111011100010100000111000100001100000100010100110100011100000000110100011111010111111100010100000001111100000000001111000001001101001100010000001101000100000000110111110100,512'b01000111111101000100000001110001110111000101010100110100111111000100110101001100110011000001110000111111001111011101010000011100011100000011010001000000110000001111000111011101000100000011110100010100110011010000000011010111010000010000111101010101110100000011001101000001111100110100110011010011000001111101001111000011010000110000110000011111010011111101000100110111010001010000111101111111001100110011010011111101110000110011111101110111110101011100010000111111010101011111111100111101011100000000011101110011,512'b00001100010000110100010011000111000011010000000100011100000000000101001101111100000000111111011111000000111101000011010000010011010100010011000101000011000011010001000111010101110001010111001100001111011111010101001101110111001101111111001100010100110011001101000000000011000100001111010011001101001100011100001101110111011100110111011100000001000000001100000000111101000111000001010011110011000000110111010100011111110001001101110001110000000101001111000101001111000101110011010001110101010100110101110001000111,512'b01000101110000000000010001000000000101000001000101000100000000110100001100001100001111000000111101010000001101000001011111001100010001001101011111000011000001000000110100111101000111000011001111110111011111001100001101011111000011110111000000000101011100111100110101001101000100010011000101010011010000111100000001110100110011000111110000110100110000000001001111110111010101000000010101110000000101110000011100000001000000110101011100010111111100010101111101010111000001110001001111000101010101000000110000110011,512'b11001100010011000000110001010000010001110000110011000111010100110001110100110100111101011100011100111111111100001100011101010001010001011100000100111101111101000111001111110011110101011101000100000000111101010011000100010111110100011100011111111101000101000100000001111100000100000000110011011111000000000001000001010001110011110100000001111101010011000100000000000000000000000001000001110001110111001101110011011101000011010011010101000000000000011101000100011111110101000100001101001101000100001111111111010101,512'b00001111000101000101000000010111111101110111110011011101000011010000110011000001011100011111000000010000001101000000000011110111001111011111000100110101011101011100111111010011000100000100011100010001000001010011000101000101010011001101111100010100110000011111001101000100000001000001010111000111000101110000110000110101000101010000000000110001010101110100001111000000110100111101000100010011001101001100111101110001010111010011110100110111000100011100000000000100111101010101111100010100010111001100110101010111,512'b01000001110111010011110101110011011101000100010011001100000000110011111101110101110000000100011100110011010111010000001101001101000111110001110100010001000011001111011100110100111101001111001100000001110101111100010111011100110000010100110000010000001111110101011111000100111101010100011101000000011111010000000000000100000000111111111100010000000000010100110111001111001111010011110100110000110011000000011111000000110100011111111111010101000101110100001100000001110101000011001100010000001101000111011111000101,512'b00011101000000010100011111111100000101000000000101000101000011110000000101000100111100011100010011011111110011010000000100011100000011000101000000000000010001011111011100011101010100010000000000010111010011000100010011110100010001111100111100111100000100010000000011010000000000010000011101000001000111010011110100110100110011001111010111110101010011011111010101111101010011000100011111110000111100000001011101001111010111011111000111110100011111010001010100110011110101111101111111010001110001111101010000001101,512'b00110111010100001111110001000001110111001101000001000101110101000000010000010100000001001100000000000001010111110011010101000011001100001101000000010100110100000101011100000101000111111111111100111100111111000001001101000001000111001101010011110011000001000011010011000001000001000111001101001100111111001100011100011100111101000101000111111111110111000011011100001101001111000011011100110100010001000000111111110000010111000000110101010000000000111100000111001101000101000111000001010100000000000000000100001100,512'b01000100000101010000111100010001110011110000110000000000000011010011000000000000000100000111000101010001000100000000010000000100011101010000000001001101001111000000001101001101110011010100010011000001111101001101010101110111010011010100111111011101011100110001110011010100001100010011010111000111111100010111000100001111111100110100010011001101010011000000000001000111001111010000000101000100111100000100010100110011010011010000000111000100110100010000111100010101111101000001111111011100111101010100111101000011,512'b11010100111111010100001111110000001111011111001100110011110000110011000000010100111101110001001100010000110000000001000100110000001111011100110100010000111111000011000100000100010001111111110001001111010000110100110001110111001101010111000100010101110011011100010000111100110101001111001100010101110111000000001100000111111111011111110011010111111101111111000001000000000000000101110111001111010000010001111100010100001100111100000101110011110001010000011111000000001111001100010111000011010101011100000100110101,512'b00011100011111011100000001001100010101010011110111000000111100000011000111000101111101000011001101000101000101001101000000110000010000000101111101111101110111010000110100010011000100110111011100000111110100010001001100110000010000110000111111110101000001000100111101110011000100000101000001001101000100110111110000001100110000010111110100011100000011010001010011110100000000001111001101110101111100000001001100110000110101110011000011110000000011010000110000010100010000011101010000001101010111010000001111010000,512'b01010111010000110001000101010111010111001111001111111111000000001100110101111100000011010000000000011111000001010100010000010000010100000001010111011101000111110101110111111100111100000000011101000000010111010101011100110101000011001111011111000001000001011111010001110000010001010011000011110100000000111100110111010000010111010000010101000111010101010100011100110111010101000101110101111111000100110000010101110111000100010001110011000000110111001100010000010011110100010100000111000111000001010001000001010001,512'b00010000010000110000110001000001111101001101010000011111010000000100111100000000111100110001000100011100001101001101010011011111011100001111001100110001001100010100010111110101001100001111110111000101001100110000111100000000011101110001110011000000000100110000001111001101110111010101110001110100111100110101010101000111110100010100110100011101000101010001000000011111110011010000011100010100001101000011110101000001011111011101001100000001010111011101000100011111010001110101010111110011000000011101011100000101,512'b11110101011100111111111101011101001101010000000011010011001100001111010111110000000000000011000011111111001100010100001111110101000011111101001101110111110001000000110100001101000100110101000011000000010101010100110000110111000100110101001101000001000111111101000000110000110000110011001101010101010111010100110001000111010100001101011111001111010011111100000011110101010101001101000111011101000001111101000101110111011101001101000001000001010001000001000000111101011101010001010101000001000100011101110100010001,512'b11111100001101000000010100010101010100010000010111111111011100110100001111000000111111111100010011110011110000001111010100110101010011011100010100110000110000110000000001001101000000110101001100000100110111001100110000111100000011000000111100001111010101110000110111110000010100000011011100000000010100000101001111110001110001000011110011000100010011110111111111110111001100000100000100001100000001001100000111110001110000000000000001111100111100110111110000110101011111000000111100010100001100010100010100000000,512'b11011100010011000011010100010111110100000111110101010101110000010101110011011101000101010011000100001100111101001100000111110100110000110111111100011111111111000001010100010001111101001100010011010000111100010011010101010100000111000011010100011101010000110001111100010100001101001111001100010011000011111101011100111101000001000101110100111101110001000001111101011100000111001111000000110001110000010011110001011101000011010001000011001100001100011100110101010100011101001100111100000000001100010001110001000101,512'b01001101010011000001010001000100000000111100010111110001010011001111011100011111001100001101011111010011010001110011010100111100111111110111111100010000000100000011010100111100011100111101011111110100001100010001000101111100000111111101001100001111011100111101010000000011011100000111001100001100000100000001000111011101010100010001010001011101011100110011110111010101111100010101000100011111001111111100110101010001000101000000111101001100000111000111011111010100111101111101000100110001111101011111111101000101,512'b01010100110011010100011100000100010111110000000001001101011100110101000000001101001111111101011101010011001100010101010000110100010111001100110101111101010000110000110101010101111101000100000000000100111100000001000100000000001111110001010011110111000011111100110100000000111101110001111101110101110001000001011101110100000111111100000000010001000101111100110000001111010101111111000000111101110111000001000001001101110011111100000011000011110011010001010001000001010011000000001111001111000000110011111111000011,512'b01000101110000011111110000011111110101000001000001110000010000110001001100010111001101111111010101000001010011011100010001000111000100010011000101110100000001011100000101111101110011000001001100011100000000000100010011110100001100001100000001010100110101010000010011001111010100001100010111011111010100111111011111000011010000010001000000110011000111000000110001110000110000111101010111010100111100000101010000110100010000110111111100111111011101010000010101000011010111010000000001010001010100001111111101110000,512'b01110100110011011111000001000100001111000001111101110101010000011101010101110100001101011101010001111100110011000000110000010100000100000000011100000100111111010111111100110111000100001111000101010001001100110011000001110011010001111111010011011111000100001100000100001100000000110001010111010011001101000111001101010100111111000111110000010101000100110011000111110101010111000111000011111100001111001100110000000000000011000011110111011100110100001100111100110100010000110000010100000111001111000000010101011101,512'b11000111011100001111010111110101001100010100110101111100111111111100110000010000000001000000000101110001010011110101110101000101110000110000111111110100110001011100111100110111010011011111000111110000111101000000000001110101000000110011011101000001110011011101010001111111111101000101001111000001001100010000010000001101000001110111111101010111000001001111110101110000000101000101010011110000000011010000110001110000011101000100001101000000000101000100000001111111001101011111110101010101110001000111010111000011,512'b01110101010101010000001101010001000111110100000011011100000000000011110001000100110001011111000011011100011100000000000011000011000100010011000011111101110000000100010101000011010001111100000001001101110000110111110000000111000011000011000000000000000011011101110100010000010111010011111101000001110011010011011101011111000100010000010111110100011101110000000101110111001101001100111111110000010001110000011101001101010100001100110011110101111100001100110111000011110101000101111100110001010000011101001111000011,512'b01010000010001011100011101111100111111011101000101000101011100000100011101010111000011011111110111001100010001111111010011110001010000000111110000011111111100010100110001001101000000010011001100000000111100011101010011110100000000000000011100011101010111000000111101001111001111110111000001110001000111110000001100001101000111001101110111000101111100111100000111000101000101001101110101110111000101001111110001000101000101111100110111110101000001110100000001010011000101110000000101001100110001111100010011000111,512'b01010011111101010101111111001111010011001100001101001100001111110101110011111100110101010011110100011111000011111100110111110100010000110100000000011100110011010000000001000000010000011111001101000001110100110100111111000100000100110001110100010001110001000100000000111100000001111101000000110001110101000100111111110100010011011111010001011101110011000111010100001111110100001100001100110100010000010011110011110100010000110100010000110111110011000011000001011111010111010011110001010111000111110011010111010111,512'b01010101110000011111010100010000000111010001010111111101110101001111010011110000011100000000110000010101001101001111010100000101110011010001001100010000011100111101110011110100110101000000010001011101010000110000000101010111110000010100010101001111110001110111010000010101000000000000010000011100010011010111000000010111000000110001000001001101010011000001001111010001000000110100010111110011111100000000001101110011011101010111110100110011110001010111000000010011011111011100000100010000111100110001111111110100,512'b01010001000011001111000100000011001111110101110101000011000111110011110000111100111101001100001111010000000100000100110000000011000111111100001100010101010001111111010000110101000101110100001100010011011100000011111100000000010001011111011111010111111100000011011100010111010000110100011100111100000000010001110101001101000000000101000001001100110011001111111101111101000001010001110101010001010011010000110011000100011111110000010101010011001100110101001100111101110011111100000111010101010000110000011100010111,512'b00010101000000011100000100010000000100000100001101010000000001011101000000111111011100111111110111010001001100000011000101110001001100110000011111000101001111000011010111001101000000011111111101000001001111000001010100110001010100010111111111000011010001011101000111010000000101110011001111111111010101110111010000011100000000110011110101010101110101111100000101000001010011111111011111001101000101000001010111000011000100001111011100010011000101000100011111011111000011001100110000000101000000000011010001010000,512'b00111101001100000100000101111100110000010000110100000001000101111111111101001101010000011100110001000101111101010100011111011100010000000001110001110100110111111101010011110011011111001111010000001101000111011100000001110100010101010101010100000001010000011101111100111101010011000001110101111100001111110000001101011100010111000100000111010001111101011100001111000001011101111101010011001111110011010011000011010001110011110100000111010100011100001111111100110111000000010011001100000101110000000101010111000100,512'b01111111010100010011111111010001010100010000001111000100000100000000001101010100110001110100111111001111110111001100110000000011001111000101111101001101001111010000000000111101000101111111001101010000011100000000110000011101110000010100110100000000010000000011010001000001110111010000000011010001110100110100010011011100000000010011111111011100011100010101001100010101010011010001000101011101110001010101000111001100110011110111010101001100000001110011011100010100001101010001010001111100010001110101000100010011,512'b00001101110000011100000100000000001100000000000011011100010100111101001101110000110001010100010001010100000111111101000101001100001111111101001100000111111111110100110011000011010001001111000001000101011111010100010111011100001100000000000001000100010000110000011100000000110011000011011101110011111101000001010100000001001100001100000000000111011101000100110101010011110111011100001111011111011111001111000011001101010001111100111101111111000011110011011101010001011111001101000001011101111100000100000000110001,512'b01000011110001111100001111001100010111011100010000000101110000110011000100110111000001000101111111000001110011011111111100111100111101110001000111000000110101010011000001000000001111111111001100000000010111110100000011010100110001001101010111010011001100110011010001010001110111010001011111000101110000010001011111001100011111111100010101000100000100010000011101000011000100110011010001110100000000000011111111001100111101110011001111010100000000011111010101000000001111000000110011110011000011110111001111111100,512'b00000011010001000111110001110011001101111100110101010100011101111111000001000000011111000100011101110001010011110000110011011111111100000101000001001111110011110101010100010100000100110001110001001100000101011100000000001100000000110101000100110111010011010100000111110000110000010001000000001111000000010000011101000101111111001100000011111111000000111100000000000111001100110000000001000000110100110001011100010100110000111101011100010100010100011101110000001111010011010001001100000011110100110100010111010011,512'b00111111111100011111000100110111110100111100001111000100000001010001000111010000000001001111000100011101000100110101000100000011000100000100010000000101001100010001000100110011110000010100010100110111111111110011001111001100010001110101110111111111110000000011110011010011110011110100010111000011001100110101010101000111010001010000010000000111001111000100000101000101010000110000111101010101010000111111010011000001000000010001111101000011010101110001000111001101010000001111001101010000010000011101000000000001,512'b00011111110101001100111111000001000001010000110100000101001100000101011111000011010100000011010011000100110100010011001111000001010111111100010001000101010111010011110100110101010000000001010101010101010011110000010000000000110001000001011101000011110101110111000111010000011111000001110000000111010000000100000000001100000011010011110001000001001101010111110100010100010111001111110111000000110011000111110001110000000011000101000011001111001100000001001111000111001100110000110101010001010111110001000000110001,512'b00111111110101110011111101001100000101011101000101000000001111000100110001001101000111010001000000111101111100110111001100000000111100001100010000111111010111111111000011000111011111001101110001110100000100110001011101010100000000010011111101111111110100110000010000110000111111111100110001110101010000000000000111000001011111110000110011001111001100010000110000010100110101110100010011010101001111000100010011010000010100011100010001111101110100000011110001000111011100000000110101010011010001111101001111011100,512'b00000101111101011101110001110000000111010000011100001111111101000011000001010001111101111100010011000000010011000100010001010001111100000011011111110100110100000000010101001101010100110001001111000011010011001101010111111100000111110000010100000100010101000000111111110011000011001111000011011100110011010000110011000111010111000100010100001101011111011101010100000111011100010011011100000001000011001101011101110011010011010000110100001111000100110100111111001101000011000011000100001100000100001100000100010101,512'b11010100000000010101111111110011000001000101110001010100001100011111000001110001110011001100000111010000110011000001010101110101110101000000000100000001110111010001000101110101110100010001110111000011010000001100000000010000110000011111010111000111000100010111110101000001110111000001000000000011001101000001000000010111000100010101000111011111110100111101110011000000110111001100111100001111010000111111110001001100011111110101011100000011111101010001010101001100000001000011111111111101010011110011010001010101,512'b01000111111101000111000100110101111100000101110000011101001100110001111101000111010100010111010011000000001100111101110100000111000100001101001100110111000101110001110101010111010011000111001100000101001111110101001111010000010111011100000101010011110000110111110111000101111100001100001101000100010100010101000011000001001100011101000111110100010011110001110000111100110000111100000000110101000011000001000000000000011111110101010100000101011100111100000000011100111100111100110011111101110011010111010001110011,512'b00000011000101110100010011111100010111000011111111000001111111010001000000001111000011110001011101011101110100011101001100000011001100001100111100110101111100110100110000000111000101001111111101000100011111110100000101000101000011000000111100111101010001111111110111000000001111001100111100110101010000011111111111110101000000000101110000110000001111001111110000000001010111111111001101001111000001010000011100111111111101000011000000011111000000000000010000111101110011010000110000000100110100110100010001111111,512'b01000001111111000100001111000111110101001101110000011101011101010001001101111100010100000011011111000111110111110011001101011100111101000000111100000011000001001100011111000000000111001111000101001101000000011111000101010101010111110011001100110011000111011111001100110101010111000111000111010000111100000000000000010000000011110100000111111101001100110001000101001111110100000100110011111100011111001111110111001111000100010100110100110100001100001111000100110111110000000000000100011101000011001100010000110001,512'b01000111111111111111110111010100000101000100000100111101000100000101000001000000110001110011000101110000000001000011000001110001000011000011010111010100111100010011000011001101010100111100110000000100001111000001001101010101110000010101000000001100110000000011110101110011111111000000000011110101000000110011110101000000110011010011001101011101110011110100001100010011110001110000000101000000000111110000000100000000010001001101010100110000010101110000001100010101110000011100011100000000000100010111001101111100,512'b01000100010011010000110000000101111111010001001100011100011100011101000000000011010000000111111101001111000000110101000100011101011101110100010111010001010101110000010011010100000100010011000100010101000011011111111111110100011111110011110101111101000001011111000101000100111101000001001100000100000100110100110000000011001101000111000000001100010000110111110111111101010100001111111111111100000001010111011100000101001101000000000111000000110000000011010001000001000100010100111111110101000011001101110100110000,512'b01110001111101110011000101111100000100010111000101110100110100000001010101010011000100010111110001000111000011000011010100010011000000011111010011110001000001000101110111011100001100011101000001011111110000010101001101001101110011110001000011010011001100011101000001111100110101111111000001110100000101111100110011000101011111010111110101011100001101000111011100010111010100010011110000001111011101010011110011011100001101111101000111000001010111001101011100110111001100000101010100010011010001000101110001010001,512'b01001101111111111111000100010000001100000101110101000101011100011111000100111100011101000000000011110000001101110111010001000111000100110111110101010011010100010011111111110111010111010111111111110001000000111101000000010111110011000000000011111111001100010000111101001100010000001100011101010011111100001111000111001111000011001101111111000100000011000100000000000011110100000111001100110111011100011111000001110000000011010011000011110001111101110001110100001101000111001111011101010000011111010000001100010011,512'b01110011000111000001001111110111001101000111010011001101001100110100000001010001000100110001111100010011000011010001000000000100011111001100111100000011011101111100000001000000111100000001111100010111110100010000010000001101000100000101110100010000000101000111110000001100001111001111001111011101001111000111111100110001010001010000000000010000010000110011110011010011001101010001110111000001110001011111000000000000010000000111010001000011001101010000011100010101110000111111010101000011001111000000010000110011,512'b01000011111111001101110100011101010111000100010000000101000001000001011101010011010100001100010100110101110100110101110001011111000101010001000101000100000011010100010101000000010001010111000100000011011100010000010101111111010001000011011111010011010101010100110100010000111100011100111101010000110101010111110000010001000011000101001100110000110101010000110111010011110011000000001111000111000000010101000001110001110100011111111100000000011100110000000011000100000000001100010101011111001101110000000001000000,512'b00000001010111010011110011111111010011110000010011010011001100000000000011001111010000001101010111110101000001110111001111001100000001001100111101010101001100010001110100110100010001001100110000001111000000110101110100000000001101011101010101010101001100010011110101111101001101000100110111001101000100010100111100001101111101010100001101010111000001011101110011111101010111000111011100000000000100111111010101010111010100001101110000010000000011010000010001000001010100011111010100000000110001001100000001110000,512'b00110000010101010111000000111101010000010111011100001111010101110001001111010111011100000000000100111100011100011100000111011101110011000100000011010100110111110100000100000101001101011111111100000001010011000011000000011100110111010111010101110000000100000001111101111100001100011100000000000001110011110100000011001100110111110111010000000000111111011111110001010011010101110111011101001101110000011111011100010011011111110111000001011111010011010001001111001100000111001111110000000101110111010000001100110100,512'b00000101110000110001110100111100001101110100001100111101110000110100111100000100000011110011000101110101000000000000000000011111010101000001000101001100111100110000110000010011110000110100110100000000000001000100111101011101000111110101111111000001000101010011110011010000010001001111010000010111001100110111001101110001001101110100111100001111010001011101001111110000000101001111111111000100000000010000010100110011001100000001010011111100111101010100011101110000001111000001010111110011001100000011010001011111,512'b11110011111111110100010111010011110000110111001101000011010000010111010100000011010100110111011111000101001100011101010001000001010011010101000111110001110100010001000111010011000000110000110011010000010001001100001100000011000001010011111101011101011111110011010011110000000111010100110101110000111101010000110000000001010100010001111111010111000111110000010101000111001100000100010101011111111100110011110011010100010011000111001100110101000001010000010000001100000111001101010000111111000000001101110011000011,512'b01110111011111000001000111001111010001110001110011010000110011010111000011110100010001000101010011000001010011111111010100011100110000000000010000111101011100110111011111011101010101010100111101000111001111000100110100011101111100000011010000001111110011110111000100111100000001110011010000110100000001000001000101110000111111000000000011001101000111110011010100010100001100000111000101001101001111110000010011010011000001000011001100001100000000110000010101110000000000110000000001010101000011010001010111010100,512'b11001101010111000001011100000011001111010011110000110100110001110011000000000000000001011100011101000111110001000101010000110011011111011111000011001100110000000111000101110101110100001101010011110000110101000011010001110101110100010101110001011101111101110011110000011101000000111101000011000100001100001100110101011100000001010001110100001101010101110100000000111101000101111101000111110111111100001101111100110011110100110001000011000000000000111111010111110000110000001100010011000000010011000100011111010001,512'b00000011011100110000011100110100010011010101111101110000000011011100001111110100000001001101010001111100111111010100011100010000000001010101001100001111001101011100001101001101011100111101110101000111010011010101000111000011000111111111110101010000010101111111000001111111110001010100010100010000001111001101010100011100000000000111000011010001001111011100110001110011010000010101000100011101000111011100001101001101010100010000001100010000000111110000000000110111001100010101000000111101000001011101010101010001,512'b00000100110100110101001100110111011101000100001111111101000001010001111111000101111111000111001100110111110100110101010000110000111111011100000000010101111101000000010000010011010111010111111111000000000100110000110001111100111101001100110111010001110100000001111111110011001100110101000011001100010100111111000101111100011101111111001101000001110101110111110111110111011101111100111111000000010000010101000001110011010000000000111111000111110101110001000011111100010000111111000100010100001100000000000001110111,512'b11000000010101011100000001000111011101011100010100110001000001000111000111010011011111110111001101000011000001000101010101110000010000111100000100010011000111010011000000011100110111000001000000000001111101110100011111001100010000110000010100000100110100001100010001010001000100011100111100000101110001010101000000000001011100010011000101000011001100010100000100011100001101001111001101110111001100110000000100000001001101000011011100111100011101010100000111111100000001110111010101110011010100000001110101000100,512'b11000111011101001101011101010011001101010011000100011111001100011100110000000011000000110101000011011101010011110111110001000000111100010011111101001100000001111100010100000011000000000100001100010011001111010111001111000011000001010001000100110001011101010001000001010011110101001111110101011100011100000101000011011111010011001111010111010011110011010001110001110011111111000100000011000100010101001101000011110000010111011100111100111111110001010101110011000001111100110111010011000011001100000100000001111100,512'b00110000000100111101111100001111011100010000010000000001000101011100010111000000010101110100110100001111010001111101111111110100110011110000000000000001010000110100010011010100010111010000010100000001010100110001010011110111010011001101011111000001000000011101000100111100110111110100010001000111000011001111000000010001011101110000000100111100000011110000110111000100000001001101010000111111111101110000110001010001000100111100001101110000000001000100001101111101110111010011011101011100110000000000010001010001,512'b01001100001100000111110011110011111111000011010100010100010001110011001100110001110011111100110101000000000111111100111101110101110100010100110101000011110101110111000000001111010001010000010000000001011101000011110101011101010101001101010000010111000101000111000101001111000111011100111100110001000000110000010000010101110100000011001101110111001111000111001111010100010011011100011111010100000111011111001101110101111101000101000011010111010101000100000111111101110100110000000111001111001101000011110111000100,512'b11001111010000010011001100110111000001010111111100000100000101000101110100010101110011010101010100110001010000001100001111111100011111111101010011110000011100110111000000000001000101111101110011001111000011000100011100010100110100001111010011010000110111111100000000111100011111000011111100110111010000110111111111110111110001110111000101010000110101001101001100011101011100000000000000111100001101011100000011110111110000000100010001001111000100110111111101110101010011001100001101001100000011011100000000010111,512'b00000000001111010101000101001101001100110101000011010100011111001100010000111111000100111101000101000100110101111101110111010101001111111100000000000100110100010101111100001100011100011111110011000100000101110000110000010101010011000001000100000000110100010101110100110100000101000000000000010111111100011101001101010100000111110101110101010111000000001100010111111101010000010000111100110011110000001100000101001101000011010001001111011111010101000111001100000101111100000100000011110011111111001111010100000100,512'b00000000000011000001010001110000010100000101010101111101011100010100000001010100111111001111011111110101010111010111000001110111000111111111000001000111110101000011010000000001011111000101001111010111110100111101000101000001111111001111000100000101111111011101110011001100111111110100000001110111000100000111110101110100000111111100000100111100000000110000011100010000000100011111111111010000010000111101110111010011110000000011001101110100110011110001110111010100010011000000001101010001110101001111010100010101,512'b11000011000001001111111101111100111111001100001111001100111111110100010111110111000100001111000100001100010011110100001101011100110100010011000001110000001111110001001101010011000101010100110100000100000000010000111111010001010101010101001100000011011100110100001100010000000111011111010100000011111101010000010000110001010111010001001100001101011101011100001101001100010100010011110001110100000001110000111100010001010001011111110000010000110011000001011111000100010000110101000111010011110111110111110111001101,512'b00011100000111011101110111010001111101001101000100110011011111001100001100000100011111010100010011010000010001010100111100000100010011000101010000000000110101010111111111001100010100111111000111011101000000110100111100001100110000001101011101110000000011111111110000010101001100110101011100111100010011011101000011111111000100001111110000110011000101010011010011000000011111001101000101010011110000000101010100000001010111010011001101010000011111000111110101111111000001000000010001110101111100001100110011000001,512'b11110101001100010011111111010101010011001101111111010111010101110111010111000001000000000001000001010000000000110001110011111100001111110001010100010100000001011101011100000101110000001111011100010001110011110000110000110001001101111111000101011101000000011100000000000001010011010111111101111100000000000100000101010011010000001100010001010101000000010001000000011111001111000001001101011100110011010101110001110011000101000001000011110000010011111111000111011101110101001111000101110000110100110000011100111111,512'b00111111110111001101000111000111110000110001011100110100111101000001111111001100110011010011110000010011110011001101001100110011000011010011110011000000010000010001111100010001010101010011000101110011010000000101000000010111010111001100000001001111110000011111110100010101111100110001010000000101010100110100000001110100000000011101111111000111011101001100010111000000010111000100001101001100010111000000010001110000000111010001000011110111001111110011000000011101000011111111000000010111000011011100010000111100,512'b11000011011111011111011100001111110101001101110100000100000001110111000011000111110100010111000111111101000000110001001100010001110000110100000000110000010011111100001101001101110001000011000111000111001111000111000101110100010111000100010000000000110000000100011100010000010111000011111100110001010000000111011101011101001101010100000011001101011101111111000001010100111101001101001111111101010100110011010101010100111101011100010101010001010111110011000001000011011111010011011100010101001111011100111111011111,512'b11110111110001110111000011110000010100000101000000011100011111000111000101110000111100000100011100110111110011000100000000000001001101010101110011110111000011110111000000110001010011000100010111001101001101010000000111001101010100000000010011010000010000001100000011010101110001110111011101111101010001110011000111111111000101011100001101010001010001000001010011111100010101000011001111000011010101110011011101110011000000001100000111010001000111000000111100010101011101011111110101110111001111010100010000010011,512'b00110111000111111111110001010001001111001111110101111100010101010111010001000001010011000000011100110100110001001100110000001100010101000000000101111100110101000000001101110001010001010001000000011100110011000001001101011101001111111100010101000101000101010000011100010111010001111100010011000000010000110001110100001111001111000100110011111111110000011100011101010011000011010111110111000101110111110011010001110000010011010000011100000101011111010111011101001111110000000100010011001111011100000001111111010100,512'b01000001110011011100111100010000000000010101111101000001110011111101000001111100110100000000110111110000010000110101110111010011111111010101111100000011000000000001001111011100110001010000010011000100110101010011001100000101001111011100010000000100000100110111011100010101110101010011000001010001000011001100000111110111000011010111010000110001001100000000000011111111111100010011000000010001111111110111010101110011010011111111000111010100110001011100010111110001000111000011010101000011000100110100000011110000,512'b01010101000000000011110111000001000111000100110101011100010001010111000011110101110101110011000001001111010011110100110001010001110101110001010000110100110000111100011111110011110111110101110000000101000000010100000000000101000001001100010011010001000111000111000001010101111100010001011101110111000001000100010100111111011100000011111101110100010111010000111100011100110100011101000001010001011100111101011101011100000101000111000000111100111101110101000011000100110011000011000000110000000000010100010000110000,512'b00111111010111111100110000111111000111110100110111110101110101111111010000110101010100110001110001110000110100111111000011010111111101001100011101010100111100111101011100011101000100000011110011010111010000110001011101001101010011000000110100110000001100111100001100010001000100111111000100110000011111011100110000110101110000000001110100000100110101010111011100010101000011001111010111111100010000000001010011110111010111000000010000000101000111111100010100001111010000001100010001111100000000110100001101110111,512'b00001100010001000100001100110001010011110011110001010000001100111101110101000001110100010011000100000100000011010100000100000101000101000011110001111100110011110000001101011100000001010011010000110101000111010011011100010011011100000100000011000101111101110101111101110001110100011111001111000101000000111101110101110100000000001100000100010011001100011100000001110101110100110000000001000101110001010100011101110001000100010100111100001100000100000011110001111100000100110000010100111100000000000101000011010000,512'b01000011010011110000010001000101001101010100001111010000000111000000000111010011000111110100110100010001000011010011001100000000001111111100010000000101000001000100011100000001000011010000000001001100011100110011111101110101000001000000110011110001010000011100011100111101000101010100011100010100110000000001111100000000011101000111110100000111000011011111000001010001001100010101000011000100000101010011000011111111010011111111010011000111110011111100010111001101000111011111000100110100011111011101001111110011,512'b11001100010100000001000000000100001111000000110111111101111100110001000001110100000100010001001111010100011101011111110001001111010100000100000000010111110000010001011111010100111101011100001100110100001101001111001100010101011100000011001100010000111101110000111111110001011100010001011101001100000011010011011100011100010101001100010101001100000100000000011101000101000011010001110000110100010000000000000101000001110011111111001111001100110000000111011101010111000000010001000000010100011111001100010100001100,512'b11000000111111011100001111110000111111111101010011110100000101110100010101001101110111110011010111110011110011000000111101001101000000011100000011001111110100110011000100110100111111110100000101001100000100011101010100111111111111110001000111111111010100011111010111111100110000111111000001001101001101011100111100111111011100001101010100000001010100111100110101000001110001010001001111000101001101110101001100010101110100110111110101110100001111001101111100010100011101110011010101000100000100011100111111010011,512'b00111101000101000000010011001101000011001111001101001111000100111101001100001101011100110011000101010000010000000100000100010011010101111101000111110011110100110000000000010111000011000100111101110101110011110011011100000000001101001111111100000000010011110011000100111101110011000011000111110001001100000000011100000101111100111111001100110011010101111100010100000101111111010111111100000101000100110000000000111111001101110101011101001111001101000001110001111100000000111101111100010011010111000111010101001100,512'b01010001110000111100010111000000011100010011111101011100010101000011001100000100000001000111000001010001110011010111001111010100011111000000001111011101000111011100010111000000111100000001000111110101010100001100010000110001110100110100111101111111000101010100110111111101011101001101110011001111001100110101001101001101110011010000010001011111011101110101010111000101110100000101000111010001010001110000011101010000110011000111010011010011110011110101110100000100010001001100010100000100011111010111000111010011,512'b01110101001100001111000111001100010011010000000101111111010100110000110100000100000000111111010100001111000000010111110000010100001100110011110000111111001111001100000000010011110111000001111101110101010000010011110000110100000011000011000111110100000011000000110000010000010101000111010101001111011101011101001111010101000111010101001100000001000000000011000001110101001101110000111100011111111111111101000111000100001100110101111111111101110011000011110001110101000000111100110001001111000011001111010100001111,512'b01000000010000111100111111001101111101011100010000110011010011110100111101111111110001010111111101010111000101010001000001000111010001011100011111111100110000001100011111010101111111000011000100110011001100001100001111010101001100011111000100111100110011000001010100000001110101000001010011110001111101000001000100000000010000000100111111000001001111001101001111000111001100011100010000110001110011010000001101111100110100000000000011010000110111001101111100000011010101000111010101011101000111001101010000110011,512'b01000001111100000111001101010000110100110000011111010011000111000001110000000100000101110011110011110000000101001101110100010000000011000100000000010000000101000011000011011100011101111111010101000000010100110000010001110001011111000100110000110011000101000001010011110111000000000011111101110011000000011111110001000000110100010011001100010000010111010111000000000001001100011111000111110101000001000001000111011100000001001111011101000101110100110100000100000000111100010100110111011111000111010001001101000000,512'b00001111000000000100110111011101001101010011110111000001110101000101111101110011111100001101000011110011000101011111111111001100111100110001110011011111001111110011001101010111110101001100000000000000011100010011111101110000110011001101110000111111011101011100110000010001000011111111000100011111010000010101111101000000000011001101010000010011010111110001000000000001010011111100000001000011010001010111011101110101110101010000110011010100000111010011001100110000000000111111010000010101010101010000110001010000,512'b11110101001101010100110011110101010001000100110101000100000101110111010100011100011111010100111100110111011101000101110100111111001100001100010011001100000011110011011111001100001101010011111100111100111111000100001100110000010000110001110100110111110011001111011101000000110011010100000011010001000000010100001100000111111100011101110011000111011111000011000001010011110011011100010011110100011111011101001100110000001100011111000011001100000100011101110000010100000000110111011111010011110000000100010001000001,512'b01110011010100110100010011011100000011110000111100001101000111111101111111111111000000000001010100000001011111111100110011111100111101010001110111111100110101000011111100000000001100011101010000010011111101110000001100110011110100010000010001110100000011010111010011000101110000001100001100110001011100000000010111110000010101001100000011000011010011000111010011110000111100011100010101000111000100010001111111010000110011010100010100001100010001000111111101000100010000010011010101110000010001001101011111010100,512'b00010000110001111101000101111111110001000101010000011111010011110011001111010000011111001101001100001101010001010100110001010111110011000000110000001101110001111101000101010001110111010100000000001101000101011111110000110001000111011111110100001100111111000100111100110100010111001111001111111111110000010011001111001100000001000111111111000000010011000100111100010000001101000001010100010111111100000001000000001101110000000011000001110101110001000100000101111100111101010100010100001111011111011111110011000111,512'b01001100010111110001010000010101000100110001110001001101011100111101010011000000000000010000010001110001010011010111011111000111111100000000110101110001110101111101110100001100110100000111110101001101000011011111010001000001010101110011110101110011010001011101001111010101001111001101111111010100011100110101011111001100000011110011010111010100010100110100110100111111000001001101010101110001010011010000110001010100010000000011001101111100011100110011001100110000111111010000111100010100000011110111011100011100,512'b00000101110100010100011111111100001101000100110001010000000111001100010000110111010000001100111100001100010001010100010000000101110100110000111101001100000001000001010011000000110100011100010000000011010101110100000111000100001101000100000001001100110101011101110000010000000100000001011101010111000100000000111111001100111101011111110001001111110100000001011111001111111101000111000101000000110000111100111111011111001111010101001111110111110100111100000100010001000000001100000001010111111100000100000100001100,512'b11010111000111111101110111010000010111110000110011000001010001010000110011010111000111000101011100001100000001000001000101010011000111110000010000010100000100010001000100111111000100010000000100010101000100110000000000000100110011010011000000011100010111111100010000111100110111110001000111110000111101010001000111001111010000000011000001000001110000000001010001001111011101011101000011110000011111010011010101011101000101000111110000011111010001110000010000010101000000110000000000110111111101001101000011000100,512'b01111111000101110011000011010111000111110000000000111101000000111101010111000100110101001111110101000001000100000111010000011100001111011100001101010001011100000001010101011101001111011111010000110101000100010000010011111111000011011101001101000000010001010100110001010000110000010100110011000101110000011100110011000111111100010100110100001100010000010100110100010000011101110101000111110111000101000000000100000000000011001101000100001111111100010101000000010011001111110000000101111100010000000001010001010001,512'b11010100110100011111010111000000010001111101000101010101111101111101010100110100000000011100110000110111010001000101110011010001000011010100011101111111111111010001010011000000000101110101000000001100000100000011000111110100010000111101010011000011000100000011111111000011000011010011001101000011010111000001001101110111000101010000010001111111000111110100010101011100000101000101001111001111011100011111111111110100000011110100010000000100110101110011000001110011010101110101110000010001010000010100001101000000,512'b01111100110011010011010011011100110000000101111100110011010111000100110000110001000000011101000001011100000001000001000101000100000101010011110011010000010111010001010011011101110001010001010100000101111100001111111111001101111111110111111100000011110101000001010011000100000011111111001111001100000001111111000001010111010000110111010111001111000101110001001111001101010000010001110111111111110101000000001111010111111111000011010011111111110000000000010000000101110111110100000101000000110011110000010100001100,512'b00011111110011010011000011000000110000110101011111110000000100110111001100110111000101011111010011011111011101110000011101001100000011010000111100010100110100000101000101110101001101110001000011110011110000001101110000110100001101110001010100011100010001000000010000111100110100000100011101110001000000110001111111000100110000110001000111010011111100010001111100000100011111000000110011010000000011110000011100010101010000011101110100111100001100110100110101011100011100011101110000110000111100011111111101000000,512'b01010001001111000000001100110111000100000101000000110101010001001100111100000011011100011111001100111101010000000111011101010011010000111100000011001111010111011101000001110001011100000011110000001111010001111111001101001101011111110100111100010101110000000000000011000011001101011111111101010101010111011101110000010000010011110001000000010001010000110000111111010111010111010000000011010000000100001111111101111111001100010111010111111100110100001111010001000100000000010100010100001100010001010101001111110101,512'b01010011110001000011000001000000111111110001110001111100011111011100000000011101010101111100111111011101110001111101000111110011000111010011000111001101000001111101111101010000010001011101110011111101000100011101010000110101111100011101110111010000011111011100110111111101110100110100110101010111011100000111110001000001010001110001010011000000000100001111001101001100010100001100110011110001000100000001000101110000110000110111111101110001110000001101001111011101011101110011000001111101001101111101001100110100,512'b11010000111111010000110100000101110100000111011111011111000101011111111100000001110001110011010001110011110101010111000000111100011111010000010001110111001101110111011101010000000011111100110011110100001101011111000001001100111100110111011101000001000100000000000100010011110111111100011111000001010011001101011100110011011100000011011101010101000101001100010101110000000111000111001101110101010001000011111101010000000100000001000100000001000011001111001111001100110111000000001100110011111111011101010011110101,512'b11001101001100001111010011110101010000010000110011010001010100010000110100110100110011001100010100111101011100011100000100011100010111000000111111011101010101001111010100111101000101110000000100110100011111000111110000000111110111111100000101010100000101010011000000010000000011000011001101010101001101110001001100011100010101010100000001001100010000111111001100000000011101010000011111000100000101110011000100000111110000110000011101010000000000110001111101110001110000001101110000110011000001110111110111000011,512'b11000111110000110000001111000100000111001101010001111111010101011111110011110001011100000100110011011111011100000111000000110001000101000100011100001111110011000000000101110000010011001111011111111101010001111100110011000101000001010011110000110111111111110000000111010101001111110011000000011101000101000100001101010011011100110011110011010011000001000001001111111111011100000001110111111100010000010000110001000101001111000000110001110011110111010011110100010100110111010101011101011111111100001101010000111100,512'b00010100000000110101110101000000110101000000110100111111010001010101010000000111000111001100110100000100000000010101010011110000110000110000000000001111000111111111000001110101011100010111010100111111010011110000010101110100001111111100011100111101110011110001110011000011010001000011110100000000000001111101010000000000000111010101110000010000000011110001110111000000010001011101000011000011111100000101000000000000110001010100011100111111000111111101000001111100010000010111111101001100110101000100000100010111,512'b00111111010101000011110100110000011111000011110000110101110000110101010011111101000000000100000011000111000001001100010001000100000000111101110101010001110001001111010100000001000111010011000001001111000111110100010001000111000111111111110000000111110001111111000011010111011100110001111111110000110101011100001100111100011100000101110011010011000001010001110001110111110001011100010100011111010100111111110111110000111100010101010011110011110101110000110000110101010011110111001101111111000101000000000100001100,512'b00011101110000110111110101011101000000000000110011110100001111111111010100000100000100010100000000110000110011000111000000000100000111000100001100010011010101000001000000000011000101000011010001010100001101110111110101110101001111111100011100010100110000001111011111011100011101000001110000000011000100110000000001110101010011011100000011110000000001001111010000111101010011001101010101010100010000010001000000111100001100110100010100001101110000111101000011000011110100011100010111111101000001011100110101111101,512'b01001101110100110011010101001100111111011111000100111100011101010011000100001101110100011100111100010011001111010100001111110100010100011100001111000000010000111100111100011100001100010000000000000001001111010001010011000111011111110100111101001101010101111111000011000001010000110101011101001101011100010011110000111111110000000001001101010000000011110001110001110100000011011111110011000001111111111101001111010011110111111101110111010001000111000001111101010011000100111100110100010011000001010001000100011100,512'b01000011010100010000110011111100000101110100001101000011011101110100000101011101000101001100000011000000000011000001010000000100001111011100110100110000110000111101010000110001001100000000110011010100000111010100010100000000000000001100110111000001110100110100010111010000110011000011110111000101111100010101000101000001110111001100010011010100110000010100011111000000111101010111000101000000000001000111110011000001001100010011001100110001111101000100011101000100111111000000011111110011000111000001001111011100,512'b11001101000111110111010000110011110100110101011111111101111101000100000000111101111100010101010101000101000011000101110000010111111100000011011100000100010000110011110000000000000001001100010000011101000001110100001100010001010011010000000000110000011111010001010000111111001100000000110011110011010001110101000111000011000011010100110100010100110111001100110011010011010011000000001100000001111101011100111111110100001111111100000100010111001111000101000111011101001111110100010111000101010011110001001100010000,512'b11010000111101010000010011000101010001001100010011110111000011000101111100000001010001111100001101110001011101000101111111001100111111000101110001010101001100111100000000010001110000011100001100110000110001000000001111110100011100000100111101000001000111000000110001110100110001000011111111110101010000001101001101001101010101001101001111010000010101011100110101010001000011010111000000111101000001010011110101010001110011001100001100001100011111110000110011001100110001000101000000000011000100010000110011110001,512'b11000100000100000001000000111100010000000100011111110000010111110011001101011100110100010101011101010000001100110111010111110001000000000111011100111101010100011101111101010000010111010001011100000011111100110000000001010111000100111100110011110001000100110000111111000011000000000011111101001101000100000011000000010111000001110000011101000001010101010100000101110001111100001101111100010101011111011100110100000101000001111111000001000111010001010011110111111101010011110001011100000011110101111111110101000000,512'b11010000001101110101011101000001001101111111010100010001001101111111000001001100110100000000011111000011000000000111010001000000010101010000110111001101110011000111110011111111010011010100110000000111001111000001000000000101010101000111110101000101010100001111000000010101110101011111110111001101000001110111001111111100001101010000111100010100010000111100011100000001010011111100010011010000110100001111011101010100110111010001000001000000110001001100000001001100110001000000111101000000010100110100000101010000,512'b00001101110001000011000100000100000100011100000101000000110011110111110000110100111111001101010011000111010111011111000101111100110000110100010111110111010111000001001101000000010100010000111100010101010100010001010101000000110011110000001101010111001100110001010000010001110011000000001100000001000011110011000001010101010100011101010000001101110101001101111111110100010101001101000100110101000000001111111101001111000100011111000100011101110100110111010101001100000000110000000011110101000101010100000000111100,512'b00010000011100010011001100000111110011110001001100110001110001000111000000111111011100010111110011110111010100110000010111111100110011000000010111111101000001011100110000001111011101001111110001001101111100000101010111110011011100110101000111000011111111010000110100001101001111110011001100001111001100110111110011000000000111110000011111110101010000111101000101010000011101000001000001000000010101000001010011010100000000111101000000011111000000001100110001011101010111000011001101110100110111000001000101110100,512'b00000100111100111101110001010000010111110100010000000111010100001100000011110111001111110111111101110011110111111101110100010000000111110101010011000001010000010000011101011111000000010101000000000100000000110101000001010111110011011100001111001111000101010000001101010111111100001101011111010100011111000001000100110001110000000100000101110100110101000000001100011111010001001101110000001100000000000011111100000001010100110000001101001101001100011101011111110100010001110000001111000000010001010101001111110000,512'b00010000010000110001010011110001111101010100110101000001010011010100000100011101011101010011010100000011000101000001110100000001110111000111010001000001110100000100110100010100110011110101000000010101110100000001000011000101110000001101110111000111011101000000000001110111110100010001011111010000110100010101011111000111110101110011111100110101000011000001111111000111110001110101011100110000000000000011110111010101000011000001000111110100010100010000011111110001001111000001110000111101000111000001010101010011,512'b11011100000011111100000101110101010000110111010011110111010101000100110000001101110101010011000111001100110001010001000100001111000111000100000000000011010111000101011111000100010001010111011111000000111111000000110100010011110101000011110100000011000101001100000101110001000000010000000000001101010011010001000000011100110101000101010000011100110100110001011101000011000011001100000101000011010000000000001101000101011111010001111100111101110100010011011101000111001100000100010000011100000001010011010100010101,512'b00111111000111000000110100000100000011000011011111011100110001010111110001000111110000110001011100000000110001110100000101110100000011010001010011110011000000010101000100110111011101011100110001110101010111010001000100011111011100010111010100000111000011000011001100110101010101001100111100011111001111010100001101110101010001010101110001000011000000110111011101110000010111000001000000000100000000110100010011110100010100001111110001000111110001001100110001010000000001110100010011110101000001010101110101001101,512'b11110001010111110000011101110000010000110100010011011111001100000111001100001100000001010011010100000001111101111111000011011100010000000011000001000001010111000011010001001111110101110100110111110011010011010111000101001101011111000000110000000001110001110001000011000111010111010111010111010111010111000101010111011101011101110111111100010000111101110001000001110101110001001100000101110100010000010000110111011101000011111101110100110101000011001111001111111111010001110100010001001111110100011111000000010101,512'b01000100011111001111000111000100110000110101010000000100110011010111010101000111110011111101110001000100000100110001001100001101000000110111010100010101110101010001110100000100000001000101010100110011001100000100000101110100010000001101000111000100110111000100010000010111011111111100010111110111000100010011110111110000111100000111000000000001010001000101000100110111010111111111011100001101111101011111010011010100010101110000011111111101001100000101000101001101110001000100111101010100110001000111010101000000,512'b11110000010111001100110101110111111101000011010000000111110001111111010100000100000000011100010011001101001111000000001111011101010111000000110001110111000011010111110111000100001101110011010000000011110000001111110011000011110000110111000001000101000001110111111101110000000001000111110000010000111101000011110001010011010001000111010000000001110111000101000111010001010001010001111111000101011100001101110000110100110000010111111101010000110100011111011101010101010000000000011101011111010000111100000101000111,512'b00010101011101111111011100001111010000110001010001110011110000110001010100010000110001001111001100001101110001011101110000000111010000010011000000110111000000011101000011110111010011000000110001000011110111110101000100110011010001010000010011001101110001111111000000001101111111010011001111111100110111111111010001110101011100011111011100000101001101000111010001001101110001000111001101110100000111000101000000000111001101011101110100001111110100010000001100000000010111010100000100000101110000000100110000110101,512'b01001100010111110101000101000100111100000001110011001111000001001101110000010001010100010101010000000100111100111111000000010000000101011100111100001101000100000100001101000000000100000100110011000000000011110000010001000001000011001111111100110011010000001101001100000011111100110011110111111100000011000100000000111100110000110000000100000000010101000000010011000111001100110101001111000101110011111100110011001100110000000101000011110000001101110011000000110111001101010011011111011101000001111101110100000000,512'b01110000011100000000110000010000001101001111001111010101000000011101011100010100110111111100011101110011110011011111010100010001011111011101000000110001011100110100110000000001111111110100110000110011110100110011010011000100000001000100010000110011110001010001000100000100110100000100000111010111110000011100010000010111000000110101000111010111000111010011010001010000010011011100000100110011000101000011010111011101010101010111010111011100001101000111010000110011001100010111010101010011000101000100011111000011,512'b00111101110000111100000011001100110111010011110001000111000011010000000111111100111101110000110101010111110100010001011111000011111101000101110011011100010101111100000001110111010011001111110000010101111111110001111111000011000011110001001111010101111111111111010011111100000001110000001111000100000100110101011101110111110011000001000111011100010011001101000011110101000101111100110011001101110001000011010101110100000001000011001100010100111100011100000101000100110111111111000111010011010000111100011111110111,512'b00000001010011000001000111001111001111010111000111001100010101111100010100110000010111110101000001110011111111111111000100001100010111110100000011010011110100000100110011010001010001000100011100010000010101010001010001110100110101000011000000110011111101110001001101111100000011000000001100110011010000010000010001000000010111010011010100001111010011011100000100001100000101110100011111010100011101000101000001000000011100111101110000011101000000010001111101000011001100001111000111001101110101110001000011001111,512'b01000101000100000111000000000001011111000001110000000000111111011111000001000111010011010000111100110011010011001111000100110000000111110101110011111100110101000011111100111111011101010101111100000000000000011100010000010011111100111100110001011111001101000011011100000100110011110001000000010000110101010101110001000101010101110011010001010101000000000000010011111111000111111100000100000011011100111101110111111100000101110000001101000000011101010001011100000001000100001111110000000100000101001100010100000000,512'b00010111001100010101110101010111010100011111111100000000110100010111110111000100110001110100110100001111110100010111110100110000000101010000011101000000000000111100111111001100010011010001011100010100110001000011000111011111110001111111110000010111010000001111000101111100111100111111111101111100010011000000000101000001001100000000000100001100010100010101010100010001010001001100110100000011011101000100001101010001000100010011010011111100010000010001001111011100001101111100011100111100000111010011001101000111,512'b11111100000001110100000100001101010001010000000000001100111111001100000000001111001100110001000011111111010100000111011100110011010111010001010001001111111111001101001101010111010000001111110000000101110011000001110101001111110011111111000100000101110101000100011100000101111100000011111100011101111111000000010000010011010001000001010111000001111100111101111101110100000011000011010001010100010111110000011101110100000001000100010001110011000000001101110111011101000000000100000000110100110011110001001111000011,512'b01000100010001000000010011110111010000010111110111000100001111000011000111000100010000001101111101000011010000010011010011110001001101111101000111000000000100010100111111000100000000110011000100110000010100000101000000110011010001110011010111010111000011000001000111001101000011110001111100011111010011110011110001010001000011111101000101111111110001110111010100011100000000000111110001001100010000000100111101011101001100001111110101000100010000110011110100010001000000000000000101010011000011110001010100000111,512'b00011100000100011111000001000111111100110011010011110000111111010111111100000100001100110000110001111101010000000011010000111111011101000111000000000101000111000011010011010000010011010101000000010001000111001111000001111101011100010001010011000000001111110011000011001111000011001100110011000001001101010001000111001111111101110000001101000000000100111100111101110000001101010100110111001101000011111111110000000000010000010011010011110111000101000001011100110000001101001101001111110001110001111100011101000111,512'b01111111000000110101111101001101111111110100011100110011011101000101000011111111010011001111010100001100110101110100001111010001010000001111000101110111110100001100110100000100000001000000000001011100110000000100000000110000010000000100011100010000010001001111001111111100110000110111011101111101001100110000010100001101000111010111010001111111110000000011110011001111000111000111110100110100010111011101011100010000000000010011010001110000110000111100001111010111000000000100110001011101000101110100110101010001,512'b00001101111111110000011100111111000000000100000100110000000100010000000101000100011100001111010100000111010001010011010101111100001111011101111111000100000100010001000001010001010000000000110100000001000101001100010000000011010100110111011101000000111111110011010011111100110100010100010111000111010001110001011111110001000011010001111101011100010111001111000101010000000100011100010100010101010100110101110011110100001111011101110101110000010001110100001111000000010100010000000101111111000001000000010001001101,512'b00110111000111001101000111010000010000110100001111000111110101110100001111000101011111110100111111111100000100111100000001111100000100010101110001010011000111110001000111110001010101010001000111000011110111010101000111010101010001110111001101010001011101011101110100110000010101111100010011000001001111000001111100110111000100010000110000000100001100110100010011010100000000000000010111001101000001010000000011011111010001000101111100001101011100010101001101111111011111000101000000011101010011111111010001001100,512'b00010000000111110001001101000001011100110011110000000100000101111101000001000111000100111101000101001100000001110001000011001111010100001111000111110101000000110101000111111101001101000011011101001100111100110001010100000000000000011100111111000011000011000000111100000001000001010111110011000001111100001101001101000100110111110100000101010000001111000011111100110001111111110100010100110100110001010101001111000100110111110000000000001101010000011101010001000100000011000001010101001100010011000011110011011100,512'b01000101011111001111010000111101111101010011001100010101000100011101001101011100010101000101001111001100111100010001110001001100110011110001000001000000000001000000000011010011000100010101010001010100010101010101000001110001000101110000010101000111000000001111001100011111011101010101110011011111010001010111010100110011001100000101000111001100010001011100001100000100111111111111110111111101110101110111110000010001111100010000110001110100110011000111011100001100010101000000001101011101111111000011010100010000,512'b11000000010000000101010001000111110111110001000100110000110101111100011100111100000001010101110001111111110100110000110100000100110100011100000011000011110001011111000101010001000000111100001111111101000000000100110001011100000001111111010011110001110001110011001111111111010001001100111100000101110111001101110000001101010001000000000100001100010000011101000000011100000001000101010011011100000111000101110111010101000101110000010011000001010111000001000101110000110000000111110011110101001101010011110101011100,512'b11000000010100011111010011110111000100110101001100010000001111011100001100010111111101010100011101010101000100110000000111110111011101000011010011111101000100011101001101110011010011011101011100000001000111110100010100001100010101000111110111001100111100011100011100110100011101110101000000000101010100110001010000000101001100110000110011000011000100011111110100110001000111010001110011000111111100110100001101110100110001010001111100000000010011000100000001001101000000010011111111000101110100010000011111001111,512'b00000101010111011101001100010100010100000000001111001111000111000011111101110100000100000111110100001101010100010000000101011100110000010001010011110111000011010100001111110100010001000000011101001101000100110100110000110011111101110011010101011101001111001111110000000000111101110101010000110000000100000000011100010100000111000000110001110001000111000100011100011101000101110100000100011111010111011111000011010101000101010011001111010011000011011101011101010111000001010001000011010111000000010100111101111111,512'b00000001001100000101001101000000010000000000010101000011110011001101110101011100111101011111010101111111010100111100011111011100111101110101001100001100111100001101000100000111111101110001110000000111010111001100010000110011011111001101010000110000001100001100110011110101000111110000000100000111000001010101010100000101000001000001110011010000111101000000000001001111110100010001110000110011110100001101110000111111011111110100110111011100011100001100010100110100010101010111000011010100110001000000011111000111,512'b01000011110000011100110000001100110101111100010011001111110111110000011111110011010100000001000001111101010001010111010000000011000111000000011101111101111101010011011100110111000111000011010000001111001101001111111100000111111101110001110000010011110000011101010011010011111100011111111100110000000000010111000000111100001101010111110101001100000111110011010011001100110100010101111111010101010101001101110000010001010011001101000100000000011100010000001100000000001101111111010011011101001101000100111101110100,512'b00000100110101110001001100010000000011011101001100011100000100000000111100001100001111110101001100011100110011010011010000111111001111000101000001001111011100010100001100010111000100010111010101111101010000000111000011001100010100000011110011001100111100110011010000011100111101000100001111011111110101110100110001010001000100110111001101000101110100000011110000000000000000001100011100010100000011010100000111000111010111001111000101010100110111010000010101000100010001110011110111111100010101000011010000000011,512'b11010101110100000000000000000100110111000000111100010011011100110000010000010111011111011111000011001111000000110011110011000001011111000001111111000011000000000100010000111100110111010000110100011100001101001100000000010000011111110111000001110001111101001101000000000100000011010100110001001100110111001111010101000011000000001100010111000100001111000001110100010100110001010101001101110001010000110101110000010011000100000100010011000000010100011101000111011100000001011100010111010011010111001101011100000111,512'b01000000000001010001110100010011010011000100000100000100110111010011110101000000011111111101110000111100111100000001111111010001000011000111110011001101110011000101000001000011000011000100010100110001000100001100001100001101010100001111110001001111011100110000000011000000000100010100110000011100110000000000110001110100010100110001110000110111110001000101110101010000010101000001111100000001110111110000010011110100000001110001011100010001010011000100010001010001111100000100010111000101010100001100010000010000,512'b01011100110000011101000000011111011101110100000101010101111101111111110100010100010111110101000000010100010001011101010000000000010100011100010001010000011101110101011101111101010011000000010111110011001111110000110011010011110100001101010001011111010001011111001101000011000011110111010000111100011101010001011101010011110111010001000101011101010001000001110101011101000100111100000011011111001100000101000100110100110001010100001111110011010101001111110001000000010001010000110000000001000111000000001100110011,512'b01010011011101010000111101110001010000000101000001111100001100011100011101000101001111111100000101010000000001011100010001000111000011110111111101000101010000110101001100000000010100000001010111000011000100111111000111001111010111000101000100110000001111010011000011001101000101110100110101010101010011111101111101111100001111000111011100000000110011010111110011001111110000011111010100011100000000000111011100000000110100000101110100001100000100000111010001000101000011110101000001010001001101000101000011110000,512'b11000000000101011101110111010100110000000111111101000001010001000100001100110000000011001111000100011100001111000001000001010001000111110000010101010011000111000100010000011101110111000000111101000001110001000001111101111111011101000000001100000111110011010100110001111111000011010011010101010000110011010111010100110111001101001101010100000001011101001111010111111111110101000100110100111111000101111100111100111101001100110100010000000011001111011100000111000011011100111111001100010000001100001101001101110011,512'b00111101000100000101001101111101010001000100000001111100011101010111000001110001000000111100000111111100110100000000110101010100011111110011001100110101000001001111111100000000000011000001110000001101010100110001110000010101111101110101111101000001000100000011010101000100110001010011001101010100011100010000010000110011000001000001110100110011110111000001110011010011001100000011110100110101110101000111001100000100010101000001000011110111011100110011000111110100111100010000011101000101010001110000110000000000,512'b11001100111111110000010100111101001101000101110100111101011111000000001101111111000011011101011111010101110101000000001101000100110000010000000111010011000111110011110101111100110100110111010000111101000001001111001101111100000011010001000000000111000000110001111111000000111111000001110001010000010101110100011101110100010001110100110100000101110101110011110011000111000001010100111101000100000000110000000000010011010100000100010100000111011100111101001101011111010000001100011111110011010111110011010011110011,512'b01000000110101001100000101000011111111000000110000110011110011110000000000010100010111000111110000000000000011110000110101110001110100011111110101010011010011000001000101111101000011001111000101011111010100000100111101000100010000010101110000001101111100110000010101110011000101111101001101001101110100010101010000000011010100000101010001010001000011111101001111110101000001000001000100000111011101110011110011110011001101000111110000011111000111010000001101001101110101010000000101001101110000010011001100110000,512'b01001101010100000101010011111101000101110001000100000101110011110101110011000100010000001111110100000001000000010100010001110000110101000011111111010100001111000011011111001100000100010000011101001100001101111101000111110000000101110000111100011111000001000011110000111101000011110001000111000100111100010000000000000100000101010111110001010011010001011100000100010000001100010111010101110000001100010111000000111100010001011100111100111101010111110001011100000111010101000100000100010011010011000000010011010100,512'b00010111110101010001000000000111000101011101110011000100001101000100000001110100010111000011111100000101001100010100111100000000110100110001110111010100110100110100110111110011000111110011010001010100010100010111011100010100110000011111010001000011000011000111111100110000010111010101010111010011000001111111010101001101011111000111011101000111110001110011011101110100010100010101111100000111000001010011010101011111000111111101011111000101010101000001000011010100001101010111000101010001010111000111001101110100,512'b01010001011101011100000100111100110111111111001101011101110001001111001111000100110001110011010100011101000001000101000000011101010011000000000101000001000011111101011101000111000001000001110000010101111100001100010000000111011111110001011101010101001111000100010011110100001100000011000100110011010000011100010111010100001100011111111111010000110100110111000001010000000001111101110000010100110101010111000001111111110000001111001100111111010111010100000011010111010111000000000011010000000000000000111100001100,512'b00000000000111011111000000000011011100001101001100010011000100110011111101111100110000000000110101110000110100010000110001001111010101000000110001010111110011000100000000000111110100011100000000010000011111110011001101110011010100000100111111111100011101000100000101000011010000110011110000010011000100000000000111110000010111110011000001110100011101010011111100000011110011010001000000011111111111110011001100010000001100010000000001010000110001010000110011010011000011000011000000111100010100110101011100001100,512'b11001111010111000100001111000000110111111101010011000001111111000000000100011101110000010011110011110011000111000001010111001111000111010000010011110001000000000100111101011111010000011101110011011101001111001101010000010101111101010000111101110111110000000111111101010001001111110111001100000001000101001101010101000011000000010001010111110011110111110111010011010100000000010111000100000111011100000111001101000101010000000001010001000111010101001100010000001101111100001100011101011100000100010111110100000011,512'b01001101110101111101000001010001000111010000110111000011000100000100010000000111000011010101000001110011110011110101000001000011110101000000111101001100111101001101010001000111111101000000000100011111001100000000010001110100011100000001110011111111111100110000010000110011000111000101111100010001011100110001110001001100110000000111011100000100110011001101000100111111000101000100000011011101011101000000010011001101110000000101001101000001110111110100010001000111000101110001110000000001110100010111010000111100,512'b01010011111111111100110001011100110100110011000011001100011111110111000111010001110111010000011100000000011111010001001101010011001100000100111100010011110100010011111101001111000011010100111111110000110111010001010011111100110000011100000000010000010101010101000011010000001101000001000101000001000001000100010011001111110100010111010011110000111111000001000011001100001100000111000000000101001100110001000100111111010000110000110011010000110000110011001100001111001101010111000111011111111100000101111101011100,512'b00000000001101010100010000010100000001110000010000000011010000000000011100111101110001010111110111011100110111010011001111000111000001011100110101001111111101000100011101110011001100110111000101001100110001010111000001110000111111110000000100111101000001001111000011000101010011001100110101110111111101111111000101010100010101010001110101000011011100000011110000010001001101010001001101000001001101001111011100000101010011000000110111011100000111110001001100000011001100011100010001000101110101110101010101000101,512'b01011101010000000111010011010101011101001100111111010111000111010001000000000000010100000000000011110000000101110011110000111100110100010001011101110001000100011101110000110000111111001111110001010111111100111101000111111111000000001100010001000101000000001100110100010011011100011101000011000100001101111111010000110001111101110011110111111111001111001101011100011100000100010011110011001111011101111100110111001111111111000101110000001100000100110011001111000011000100010100111100000111000001010011010100110011,512'b00000011010100000000111100000011010000010000110000000001000000010001010001110011001100011100010001000100000000000100000000110001011100011111110101000111001111010101000011000111000101000111000111110001000000010011001100110111000011010001010000001101110011110001110100111101111101000011111101000011001101001100010111000111000000110011010001110101000101110111000001000011011100010100111111010101110001010000000000000111011101010000000111110111001101000000110111110111110100010101000011110011001100010011111111111111,512'b01110101001111010001001100111100011101110011010111010100010100110111011111110000000100111111111101010000000100111100001111000000000011110100010101000101011100010000010100010001001100111100010101000100111101000000010101010111110101001111110001010001111100000000010100110000000100010011010000111111000100000001111111111111110001000101010000010000110100011111110101011101000100000011110111110100000011000100000100111100001101110000001101011111000101010011001100010000000011000100000011110000000100001101110011110111,512'b00110000111100110100110001011101010011000111011101010011110111001111000111000001110000000100010000111101000101010000010011111101110100000111001100010111000011111100010000010101010111010001001111111111000101111111010000110111000011110000000111010011001101010000000100111101001100010011000100001101110000000011000100000000110001111100010100111111001111110001011111110001011100001100010100110111000101001100011100010100011111011111000111110000110111010000110011010001001100010111011111001100000000000101010111001111,512'b00011101111101011101001111010000000001010011001101000101110011010011110111010001011101000100001100000011010111010100000111000100001111011100011100000001001101010011000000110011110100010100001111110111000000111100110001110111010100001101001100000100001100010111110111110000110000001111010001001101110111000100010000000100010011010001111100001111001100000011010001010011000101110111010100000011000011110000010111001111110000111111000100111101010101011101010111000100010100000101001101110000001101001100000100000100,512'b11010000011101000111000000010100001111110111110101010001000101011101011100110000001111010011111101010001011101110001011101110111011100010011011111011111110101111100011111110000010100000000111111010011001100110111010011011101001100010100011100110000110100001100001101000111000011110001010011110101000001000101010011110111000111111100000011110111000111000011000000011111111100111100110000000001011101001101110001010011011111010101111101110100110000000101000011111100111100010001000000110011000101010000000011010011,512'b01001100000001001101010111110000010111000111000100110000001101110100010000011100011111010100000011000101110001000100110000001101000100010001110101001101110000010100010111000101000001001111010000110111011101000101111100110100011101000111000111010111000100010100000011010001001111010001011111111111001101110100111111110011010100111100000011001111111100001100000000010011001101010011111100000111001111010100111100111100000011111100111111010001110011010000110101001111011100110111000000011101111111010100010000111100,512'b01110000110111110111011111010100111101010100010000000000000101000011110011001101000100000000001100000100110011011100110011010011010111000000000000000011110000110001001100010000000111000000001111010111000001001111111100000101110001010111001101111100000011110000010000010001001100001111010011000100010100011101110000110101010011001101001100110000111111110011111100010111110111000001000001000101000001111101010011111101110111000101000101010000110000000001010101110001001101010100000011011111001111110111110101010111,512'b00011101010001010100010000000101000000111111110100000111011101110111011111110001010011110000010101010111010101010011110001000101000101000111001101001101001100010011000001011101010000001111000101001100110101110011111100010001111101000111010100010101000111010000110000010001110101001111000011110011010000010001000000001101001111001111001101010101010000011100000011011100010111000101010111000111000100010101000001011111111101000111010000111111000100000101010000111101000011000001000100000011000000011111001111000000,512'b11111100000011000011110011111111001101111111000111111100001111000001001111001100010111111100010000110000010101000111010100011101000000110001110001010000001101010000000000000001001100000111010000111101000000000000010011010101010001011100000000000001111100010001000000010000011111110100111100001101010100110101000100011100010001011101001100000011110000000111110000111111010011011100110000000100011111111101110000000101110001011111000100010000001101110100010100010100110011111101111101000000110101010011110100111111,512'b01010001110100011100000000000001111111110111000101010000110001010101000111111111110000000000111100011111000111000011111100000001110000110101001100000011110011001111000100011100000000001111010011000000110001010000000001010111110001001100010000001100001111001101110001110000110000111111010001000001010101011100010000110100110011111100011111110100010101011101010000000011011100011111111100110001110001001101010011111111001100001100110111001101110011010000110111000011000000010101011111000000000100010101000000000100,512'b00000101110011010101001111000101011100001101001111110100001111000101010011011100000100010011001111001101011100000000010111000011001101011100110000011101011111110000110101000101000001110111010111001111010000010100000000010111011101000011010000111101110100011100001101000000110100010011000000110000000111111101110100110111000101110100110100110011010111110011110111000100001101000011110000110011110001110101010001110100010100000011010101000001001101111100000000001101010100000000000011000000000100110001000001111101,512'b00010100111100011100010001001101001101010101010000000101000011010100000001010001110000000000000000010001000011000000000001010001111101001111010000110111111100010011111111011101001111111111001100001111000011110101011100010100000011011100001101000000001111000101110001001100010001110011111101000001011100011101011111110100010101010001000000001100110000111111010100110000110111110111010100111101000100000011001111111111001101001101010011110011010000110001010000000000110001001101110101000111010111010001110100011101,512'b01110101110101000001000101111100110000001101011100000100010000110001000011001100011101000111010011010101001111011101110100010101000000000000000000010111001101110011110111110101110111011111000001011111000000110101110101001101001100010111110100110000001101111111110000010100010111110011010100000000110101000000110011010001001111000111001111010011111101000001000101110100110000010001011100110101000000000100000100000101000011010101011100000111010001000101000011000011010000000011110111110011110100010111110011111100,512'b00000011001100000111010100111101001101010001000000111111000000110100001100110001010000000000010111110011001101110000110111010101111101011100000000110111111111011111011111011100110101000101110100110111110101000011011111110011000101001101001111000000010001010001010111001100010011000000000100001100000111111101110001001100111101110011010000000001010000000111111101010100110101000111010101010000000101010100000011001100000111000100000111110000010111011101010100001101011101000001110100011100111101110111001111000000,512'b00011101111100111100000000000000010100000111010011111111000011110100000100000011010100001100010000110000010101110101110000010101110001001101011100111111000011110100011100110011000101110100000111010000000001011100000000000011110000110111110101001100110101011100000100010111110100111101110011000111010011010011111101110101011101111100010101010111000101011101110001001111010101010011010000000101000100001100111111000101110111010001110100010011000011010100010001011101110100000000000101111111010011011100011100110001,512'b01001100010111111100110001000111110011000001010000000000010001010111000001110000110111111111010001010111111100000001010100010011000011000000111100001111110101000001001100010001111101110111000011010101110011110011010101001100001100000101010001110100000111000001000101110111010111010000000111010100011100011111000011001101000001110001001101110001000101001100110011000101111100001100001100010100110011010100011101000011001100110011110011111100000101110100000100111100000100010100110111110100010011110111011100001101,512'b11001101010101000000001111111101011101110101010011000000111111110000011111000001011101111111011100011111110011000011000111110100111111110101000001000011001101000000111100110011110100000011110001010011001100110101001100110100001101000000000000011111000111011101011111001111110011010000001100111100011101001100001111110111000111011100000000011100011111111100111101000000000111000001010001110011111100000111110001110101111101000100010100110101001111110011000111000101001100110000011100010000010100001101010111011101,512'b01001111000100010101111101001100110001010100000011011100111100010111010101001100000101110000000100111111000000000100000101110001011100110101000100000011010001000000000001000011110000000111011100000100010000010100110000010011001101000100011100010101110101010000011100010101111101111100000101011100000000110111010011011101010101010000000100000011110111010000000000010111110111000100000001010000110001111100010000000000010100111111010001001101000111000001000101110111001101011100001111001101000001111111110001110100,512'b01010100110111111111000001010101000100001111011111010101001111110111000001000001010000110001010100000100010111010111110001000001111100011100010000001100010101111101000011001111010101110000010100010001011101000100000100000001110001010000110011011101110000110101000000110100111101000000010001000111000001010111010111110101001111000000011111010000000011111111001101000111000100010101110100010011110000001101000111010111001111111101000000011100000111010011110011110000010000010001110111000011000101110001001100000000,512'b01001100110001000100010011000011110111000000110011010011111111001111110000000111010000000111111101110100000001000011000100011111110011010000010001010001001101000100001100001101000101010000011111110001011100000000110101001111000100110100010100011111111100000111010000110100000001110000000101010001000000000011010011000111000100110001111101110011110011010000110000000001110001001111000001011100000000011101110101110111010011001101000000010111000101111100010000011100000111011100110011010111000000110011000100000101,512'b00110000010000010111010100010100001101000100110100110101011100110100000100000001110000010011000111110101000111001100000011000100111100001100111111010111111111000000001111010100110111001100111111011101010111001111110000111111000101110101010011110101000101010111010111110001111100010011001101110000110011110100011100001100111111010111010001010100010111110000010011010100001111111111010000011101110111111101000001001100011101110001011100010111000111001111000100001111000100010111110101111100110100011100010011110100,512'b00110100000000010100000111011101110001001101001100010100011100011100011111001111010011000111000000000000111101110001010011001101010011110011010001000011001111010100010011011111011111110111110101110001001101000000010111110011000011000100000111010001001100110100110101010000001100001101000000111101000111000111000011010000001101000100011100010111000111011100000011010111010011001111000111000011000001111101000001000100010101000001111101000100010001010000001100110101111101111111010011001111011101000100011111011101,512'b11010011001100001111010101000101001111110000110000011100010000010001110000001100111101110001010111000000001101010011011111000000010111110001011101011111000111011100010000110001111111000100111100000011111101010101000111011100110011110111010101010111000111110101010101010000010001011100010011011101110000000111110000111101010011111111111101110000000001110101001101010100001111000101110001011101000001110000011111001101000000000101010001000100001100110100011100010011110100000101011100110101000011110011010100111111,512'b00010100011100011111001100000101000100010000010001010101011111010011110101110100110101110000000100011100110101000001001100001101000111000011000111010100000000001100001111110100011100011101001100010100110000000011110000000100000101000011001111111111110001111101000000010001000011110111110111000000010011110000000011000111000001010101000101110111110111000100011111000000001100000011000000010111110000111101001100000101000001001101011111110011110000001101000000010111000111000100110100000000011111000101110101110011,512'b00010001010011110011001100111101110111011100110111010000010111000100000001010100000100000001000001000111000111110000000111010011111100111111000001111101000011010111011111010000000011000100011100000001000001110101010111010100000011010011010101110101110011010001110000001100110000011101111100000000111101001111001101001100001111110000011111111100000000000101011101000011001100001100000001010001010111011100001101110111000001000101010011110100010111000011000101110001010000110000011100000011000100010000000000010101,512'b11001101001100001101000100010100111101110100010100000001000011000111010101001100000001110001010101000000011101010100110011011101011100000000000011110100001101001111010111110111000101110101011101110000011111110101000111010111111111011100110001001100110000110101000100011100110000010111110011000001000011010100001101011111110000111101010011110111001100110011110100011100010101000001000111110101110001001100110111110000000000010100010001000100110000000001111100000001111111110101110100111100110000000000001101111101,512'b11000011001101011100001111110000011111110000000100110001111111010011011101000000010100000011110000010101001101110001000001111111111111000001110000111101010011111100000101011100111111000001010000000001001111000101110100111111010101110011110111000000110011111100010001001100111111010101010011110000111101000001111100010100110101000100011111010001000000001100000001001100011100000001110011111100000000010100000100110000000000110011000011011100010111111111010011010000000000110101010000000100001100000000010001000011,512'b00011101111100110000001111000000000011010001010011010111010101000101110011001100010011010111011111110000011111000000001111010100001100111101110000110001010100010011011111000011010100010001011111110100000011010100000001000101011101000001000101011100111100000000110100110011000000000001000011000100010011000001110100011101001101000000010011000101110101001101010111000000001111000100110101000101001101001111000011011101010001111100111100001101110101110001011101010011011100000100010100000000000101110000000011110011,512'b01110000111111110001001100010000111111010100000000001100111101011100010100111100000001110101000101000101010000010011110101000100110011110101000100010101110101000001010011000000010001010100010011010111000011000011110011001111000101011111001101010000010000010001000111011111001101010100110100001100010011110100110011111100001101110011000001010101110000010111110100110111000011011111110101010001000100011100000001000011000101110001000101001101111101000101110111111100010101110000000000001111110011000011010100001100,512'b11110000010011000100000100000111010101000100110111010101111111111111000101010101000011010011010000111101000111001100110100011111011101110011001101010001111101001111111100001101111111110011000100010000000100110100000001011100110101000001000111011100010111010111110101010000000001000011011111000100010000110001110011000001110011000111010111000001011111010111001101010000010001111101010111001100010011001111000001000000110111010001111101010011110101111101011100000101010100011100011100010011000101010111011111001101,512'b00110101010000010111000001001100110011010000000111011111111111110100110000111111110101010100010101001111000011011100000100111111010001011101000011011101001111010101110101110000000001000011001101111100110000001111000000010111111100111101111111010101010001011111011100010011011101111101001111001101110100000000000101000000011100010000001101111100000001110011110000111101111101010101010000000001110100000100011101000100000101001111010011111100011100000011111111010101000001111111000111111101110111001111000001010100,512'b01110000001100000111001111000100010100110100010001111101110011001111010100001111110101010001001100010100110001000011010000110101110011000001000001001100110000111111010011000000110100010001110111110011010001111100010000011101000000010101010100000000110000000101111111001101000000000101001111110100000001000100010000000001001100000111000101011101000111110101110101010000010100010101000111000000000000110000000101000000011100011111001101000111010101000000001101000111010000001101010000000101010111010101001101110011,512'b11000011110011011100000000000101011101001100000001110000001111110100000000000100010011111100011100010001000100111101011101110111000001011100110000000111001111000000000011010100110111110000000101110000000000000001010001000001000101010011000101001101000111110111010001110001000001000101011100111101110100001111010001110101011100000001000111000111110001010011010100111100000011110111000011110000011100111101010100110111001101000100010001011101010100110001010011010101011100111100010001000011010001010000110000110001,512'b11001100010001010001000000011100110111000111111101111101111111110011000011000001110101000101000111000000110001001101110000011100110000001101000000110101010101110101110111110111000011001100010001111111111100010111000011010000000000111100000001010000111111010001010011001111001111110100010000000001000100001101010001000000011100110000000001000001111111000001110100010001010011011101000001000111000101110000110111000111000001001111000101011100010000110001110111010100110000111101110111011111000000010001000001000111,512'b01110100010001111111001100001100000000110000000011111111011101000111000001000100110011000101000001000100000011000111110000110100000100001101010100110000110101110001110011011101010100011100110111111101011100010011000001000101110011111100110101011101011101001101111100000011110011000100010100010011010011000000000111001111010000000101111100000011000000110011001100111111000001110111000000000111010100000000110000110101011111110011010111000000111111000001110011010001111100000100111111000111001100001101110001010000,512'b01011101000111001100000001110100110100001111110101110000011111001111010001000100000101010100000000011100001111000100000100011111110101110000110100000101001111010101011111110011000011000001010000010100110011001100000100000111000100010000010011010001110001000000001100000111011100110000110001110000001111010011011100001100011101010011000100110101010100010000010000000000000111110011110111011111000001110000000000001100010011001100010111000101000100001100010011010111000100010111000011010011001100001101010001000011,512'b00110100000000010000000100010100000001011101010011001100110000110111011111110011010000001100000111111100001101010100011111000001011100001100000111110000111100010000110011000111110000001111000000010101000001110011010101001100000011000001000011000101111111000100000011000100010111001111010101000100000001000000010101000000001111011111010000001100111100011111110100110000110101010011010011000101111100001111001111011100111100110011001101111111011111000101011100000101011101010111110111011111010000000100000000000011,512'b11000101000011010111110101000011011111000101111100010001000101000100000111001111001111001111000011001101010100000100001100000011010001010101001100000011010001110000110001110111001100010000111111010011000001010011111100110011010000110001010001000011000100001100000001110001010000010111000011011101010011111100111111110100000100010001001101011100110000000100000000001111010111000100001100111100110100110101001100000001001111110000000001000111110011111100000100010101010001000000011100111101000001000000111101001101,512'b11000000000000000101000011000001011111000111110011110111000001011111110000010111110000001111110011000001000100111101010001001111010101011100111101111111010011110101001101011111000100011100000101011100010000011100000111001100110111011100000001000100001111110001010101011101110011111100010011001100000001010101110101110001000111111101110100000001001111110111111101110000000011000111000011111111111101110001000011111111110000001111010100111111010011110011000100000101110101110100111100011100001100000100111111110111,512'b01011100110100110100111101001111010100000111010111111101001111000100010111000011011100011101110101111101011101110111110100011100110011111101000011001111000111001101110100010011010011000000000101000011110111111111000000111101111101010001010000010101000001110100001111000101000000110001110001110100010000000000000100001111010001001101110101000001111100110001110011010001110011000100001111011111000111010101000000000000001100010100000101111111001101111111011100001111000000000111110100001100010001110000110011010011,512'b00110100000011111101010111111100111100011111110111001101110000000111011100111101010100001111000001010111010001111101000111010001111100111101010001011100001101010011110100001111011100000111011101001111110001110000010001000101000111001101000100110000010011110100000101001100011100000011000011010001001100010011011111010000001101011100000100011111000100011111110000000001001101000101011100110101011101111101001101001101010000000100011100010001001101010101011101110000011101000100000000001100011101010000000101000101,512'b11010101000100110101110011111100010001110001000000010100010111001100001101000111110000000011110100110100000000010011000101000101110011000001001111001101010011000101111101000011011101011100111100110111000001010111010100110011110000000000110111110101011111000111010001110011110111010000110000111101111101011111010111010011000001110101011100110101000000010001000100001111010100010100010100110100110111000000000100110000010101111101111111110000111111010111010000010001010101110001010101001100010001011101000011010000,512'b01000001010111111111111100111101001100010000110001010111000001111111111111010100010011110011111101010011010000000101110000110100011101111100001101110101010001001111110001110000110001000100110000011101110100110001010111000001110001110011011101001111010100001111000000010111110111111111010101110111000100110101000100010000001111001100010100011111000001110011110011010001010000110101111100000001000100110111010000110000000100111111011101110000000011110101110000000001011111000100001101000100000111010000001100000100,512'b00010100110001000001110101011111000000000111010100110000010000000001110000000011011101110001010000110011010111111100010100110000111111110011110001001111011101000000110111110100011101011101110111000000000000000001011101111111010000000100110101011101001100110011110101000100110101010111011111010111011101110000110000001111000000110000001101001111010001010101000011001111011100111100110111000111001100001101110100000011010000011101111111110000010001110000010111010000011100011100010000000111110011110001111100111100,512'b01010000000001110001001101010101001111010101110000000101010011001101001111011111000000111101000101000101110101011101010101010100000011010011010100010111000011010001110100011101011101011101111100110000000011110100110000111101110001110101110001010000000111001101011100010100001101011100010100110100000011000111010100001100000000000100000001010001011101110011011101000000011100011111111111001100010001000011010000110011110001011111111100010000010100000000000001000000111101010111111100110011110011000100010111011101,512'b01011101010011000011001111111111110100110100111100110011000011000011000011000111010001110011001100111100000000000001011100000000010000000001001101110000110000110101010100010100110011110000000101110101010100110000010011110000010000011101000000010100001100000011010111000011001101010100000011011111000111000001111111001111110001000011000000010111011101000001011101010011001101000111010111110000010101001111110000110011110001011100000100011100110100011100010001110001001100010001110001010111110011010100000001010100,512'b00110000000100010101110011111101010111001101110000001100000000001100111101000000000011011100000100010111000011111111001111011100000101001111000101010000000111110011110000010101110000000101000101000111001101010000110011000001110000011101110011001101001100110100010111001100001111011100011100110100001111010100001101000111010000000011010001000101010111000000011101001111011111111101010001010000110100001111001111000111000100001101111111001101110100000011110100010111000101111100111100010000000000001100110101000111,512'b00001101001100001111011101000111000001011101000001000101000000110011010111000011001101010101001111000011000001010011110100110100000111110001001111011100110100010000110000001100001100000101010111000100000100000101001111110011010011010001010101001100111101000101000001010111010011011101001111001111001101000011010101110011000011110000000111110000000000000111010100110101011111010100011111001101000001010000000100010101000001110100110001000100001100110101111101010000110000010001011100011100001100110000000111111111,512'b00000000110000010001010011010111011100110111111100001100010001111100110011000100000000011101010000011101011100010111110101011111000001111100110000011101010011000001010100010101111100111111000001110111001100010011010011011111010011001111010000110100001100110000010100010100001100000000000011010001110100010111011100000011000100110001000000110100000000011111010100110001000100111100010100001100000100010101010011011100000001010100110000001101110101010101011100110011110011111101010000010111000100010111000001110000,512'b00000100010100000000111111010101010001000111110011110001010000110100011100000000110111000000011100111100110000111101000000110100000100010100110101010101001100010101110011001111110100001101000100110011110001010011001101010100110101011111001101000000010111000001010000111100010011011111000011010001110101001101010001110100010000010111000001011111010011010001011101011100111111010101111111010101110000010001000100110101010011010111110101011100010001000100000101000001011100000111010000001111001100000101110001000001,512'b00110000010000111100000100000101011100000111010000011101011100001101001100010111110101000100110000010100110011111100000001011100000011110011010000110011110101001101000101111100000100110000001111110000011100000000000011110101011101010101110100110101000101001101110101000011010011000001110101111101110111001111000001001101001101011101111111110100000001000000110011110001010000010000111111010000110011001101011101111100000011011111111100000101001111110011001111010111010100001101111100000001010101000001110011011101,512'b11111101000001001100010000011100000001001101000000000000011101000100000001001101010001000100001100010000000001010000110001010101000000110001000101011100110111000001110011010111001101011111000011000011010001011101110111110011010101000011010100111111110100110100001101011101010101011101000000110000010001110011111100010001001101000011000001010101010000011111000000011111000000111101000000011100110011010011010011001101111100000101010000001100010000000000010100011111000101000001111101010011000001010011010100010011,512'b00010001010000010001000000110101010001110100000000000011010000110001000100011111010111110011000011000001010011110100000101000001111100010111011100000000010011000011110100110111000101010101011100000011001101000011010100000011111100000100000011111100000000011111110011001100010001001101001100000101110000000101000100111111000001111111110100001100010000011111111111001101111101000111000111111111110001001100010101001101111101010011110100000111111111110011000011010101010100001111000100000111001111110100000100010001,512'b11010001001100110100110000000101111101010101110000010011000111000111001111000100010011110001110000110111010011010001111100001101010001000101000001000100000111000011001111110001000101001111001101011111010011000001011101010101111101000000001100110100111111011101000111010111110000110001110011110100000000010111010001001101000100011100010101111101110100110011110100010001010011011100010100010111110111110000000000110100010000000000111101110001110011011111110011110000110000011101010001110000000001110001011101111101,512'b11111100000100011101110111000000011100110000110101011101011100000001011100000011011100011101110000001100000100110001011111111111010111001111000100001101011111010100001111111101011100000100011100110001000011000100000100010100000011011101110000110111110111010111110011000111000011000101010001000100001100011100001101000011000001000011111100111100010101011111001101001100000100110000011111000000000101110100010001110111001111110000010000111111010101010100110100011101001111000011000001000111000101010000000000000101,512'b01010011001111001101010101001101011101010011000100110111000000111111110000110011000000010100011100000111111100000100000001110000000011010101010100010111010101110100110000011100000011111100110000001111010011001101000000010001110000110101000001000111010111010001000101110100010101111100000001011101011100000100001101111111001100010000010011110011010011000001110101010111000101000001000001010000111100010001111101010101000001010111000001010100001100001100001100000001001111111111111111010000000101010001000000111101,512'b01001100001101000111111100010001000000010100010000111101011111010101010111000011110111110101011101000100000000001100110000010100111100010100000101000111011100110101110111001111111100110000000011000001110001110101111100000111000000010001000000010100000001010011001111110001000000000001001101000111110001110011000011000000010000110000010100010100000001111111111100111100000011000000111100110111001101110100001101010101000101010000000111000011111100001101110011110111011101110000110101111111111101010111000001010001,512'b00010100110000010101010100000111110000010111000011110000110000010001110101001101011111000001000100000011000101001111010011011100000000010001110100110100001111110100011101010001110000000000110111110000011111000001000100001111010011000111010100111101010101001100111100000100010111110011010100110001010001000000010100110000111111110101000001110101000011001111000000000000011100011101001111110111010001110100110011110000000001010101011101111111000001010111011111111100001100001101001111111111111100010001000001001100,512'b11000100010101000000010111110111010011010000001101111100011100110011011100110000011100010100110100110011010111010001011101000001111111011100001100011111010011010111110001111111110011110001001101010101000000111111000011111100111100000111011101011111010001111101110100111101000100001101110001110001000011111111000000011100001111001101110011001100000100001111011100011100010101010101110011000011010000010000010011111100110001000111110001111111010111001100010000111111011101010011111100000001110111010111010001001111,512'b11010100110101110000001101110101001101010101000100000000111111000000011100110111111101110011110001000111110000110100000111110100111100110111110000010100010111000001001100000001010100011100010101001111110000010100110111000000010111010011110000000111001101010011000000011111110101110101000111001111000111111111011100010100001111000001010000010111010000011101000001000100111101011100110001110100001111010011001101010111010000110011110001001111111111001101001101000100011111001101000111111101010000000000110111001100,512'b00000101001111110000111111010011110100000011010000110100000011110100000011010111000000011111000011110111011100010100010101000101110000000000001101010001110011111100000101001111001111000101110100110101000100001101000100000001000100010101000111010000011100110101110101000011011101000111111111010001001101001100010001110101010111010111000001000111001100111100111111000101000100000111000111001111110111110101111111000111000011110011110111011101110011010000010011110100110111001101011100001100010101111100010001111111,512'b01111100110101110011000100001101110011011111001100110001000100011101110111010001010101001100010000011100111111110100111100000001111101010011001100001100001101010111011100010111011100000001110111010000000100000100010001010001000000010000110000110011000101110001001101111100001111110100110000111111011111110111110011000000110000010111001100000001111100111111110100110000000000010001111111000000010100001101011100010100000100110011111100000000110100010001000001111100111100000000111100000011111111000001011100000001,512'b00110000011101010100000000111100111101000100110011001101000000000001011111111111110001010011011101001100000111000000000000011111000000110000010001111101010101010001110111010101010101010001000011010001000000010000010111111101111100000100000011000011001101000011000000010011010111110111011100011101110001010111111101000000000000111111110001001111000111111100110000000000011100010000000001010000010101010111000100001100010111010100010011111111000100111101010100110111001100110011000100000001000111000011001100110000,512'b00111100110000000100001101110001010011111100110111001111110111011111000001001100110100111101011101010000011111000101000011000011110111110101010000110000110001110000010001110101010000011111001100111100010001000111111111000111111101111101110100000111110101010101110100000101000001001100010100010100011100000000110011110101011101010011010100110100110101010000011101001100001111110011001111001111110100010100000011110100110001110000001100001101110000110101111111001111000111011101001111000001110011110011110000010000,512'b11110001111111110000111111010000000011000000110100010111000001110100010101110100001111110100110101000001000100000100010111000100001100010011000000110000001111000100110000010011000100110111011111000111010001000001110000110000000000110001010000001101000001110011010000110100010011010001000001010100010101010001000111010100110001000000001101001100000011000111010000000100110111000100000101111111000000010000011101110001110001111100110011110100010100111100000101000011001101010001011101001100000101000011000000011101,512'b00001100000101001100010101001111000001010001000000001111011100000101000111000111110111000001010001110111110000110101111111011101000000000011010011010101110111110101001101000101110001110001010011000011010101010011111100110111000101000001110111000000111101000001011100010000010000011101000100010000010001011101111100011100000001010001000011001111110000110000000000011100000101000001000101000101010111001111000101000011000001000001010100000000010011000100110000010001111101000101000101011111000011010000001111011101,512'b00010101000000011101000001010101110011110011000111110100010000000100110101001100111100010000011111110101011111001100011100001111000111010000001101010000111111000000000000000101000111010100111101001111001111110000010101111101000101110100001100001100110111000111000011110000111100010000010100010100000111000100010111000100000100000100000001000000000011001100010001000000110111110001000101001100110001110101010100000100000111110000000000001100010001110001010101111100010111011100110111111111010111110000010011001100,512'b11001100110101001100001100010011110000010101000001110111110111010100000000000111000101110100001101111100010011111100011111010001010111110011111100110000111100000000011100110000001100111101111100111111110100110000110100111101110101011100000100000000111111000011011100110000001100000111010001010011010001001101010001001111000111010001010111110101010100010000111100000111110111011100001111001100010000000000111101010101000101000111001101011101000111110111110101000011110000001101110011110000001100001100010111000111,512'b00000001110100010011010000000001010001000011000111000011011101111111110101010000000111110011010111110000010000000001000101001111110101110111010000011100010001111100000101110001000011010000001111110001110001010000000011111111110100110011011100110000001101001100000100001100110001010100110011011100011111111100110001110100000101010000000111001100111101110011000001011111000101111100010001001111110011000001110000110000000101000001110100000101110011000111010001110011110001000101001100110001110011111111011100110111,512'b00010011000011110100110000000111000100110101011100001100110001001101111111010101000101000001001100111111000000110000111100110000000001010101010100001101110111110011011111111100010011110011110011001100011100110011001100010000001101010000110000011100010001110100011101111101110001110001010100001101011111110000110000000000000100111100000000110011011100000111001111001100111111110101011100011111001100000001110001000111000101001101110101011111011111000001000100010011010111001101011111010001111100110100110011000101,512'b11011100110011000100110001010001010011111111110100001111110101010101000001110111110000110000110001001111110011010000001100010011010101000001110000110001110111000100010100010011110011110000111100001111110000110000110001110100110011111100000111110000000011000100000001011111010100111100110111110001011111111111000011001111001100010100110100000100110000010111110001001111000001000000000001110101111100111111001101010101110011010100010100000101000011000101000001010101111111010000010100110100110011000101110011110100,512'b11000111110111000100011111110001010000110001010000110001001101000111000111011111010111110011111100000000010111001101110100010011000101110101010111000011010000110101000111010001000101110000111100000111010101000000011111011101001101000011000000000101110100110001011100110101001111110000000001000000010000110000000100110011110101000001010011010100111100111111110011011101110011110101001100000011000000000101000000110001000101110101000000000000000011011100001100010111010011110100111101000111001100110011010100010011,512'b00000100001111110111110000000011110001011101010101001100111101111111000101000011000001111100000100000001111111111111011100111101111100110001010100110011111100111100110001000001010011000001010100011111110100110111111100010100000000110100010100110101111101000100111111001111000001000011110000111111010000001101010001000011010101000001000111010001010000010011001101010000111101110001000000111100110101000001111101110100011100110001001100000111110001010011000101110011010001110100000101011111011100111101001101110001,512'b01111101110000001111110001011100010101110101010000010100001101010101010111110100110100010001000001110011000100001111000100010111000001000000110111011101110000111111010001010111001101011101000011010001010001010011010100111100011111010011110011000011111111110000111111010100110111000100001101000111010001110011001111011100011100110111000011001111010100010000010111000111011100011100010001110001001101010011000001010100110101110101000000000011011100110000110000010001010001111111111100010011110011111111000011000000,512'b11110101010101010101010000011101010101110100010111001111111100001111010001110001000111110100000000110111001111110100010100010000001100011100110111010000111100001100110111010011011100111101011111110001000000000001110100111101111111110011001100110011010000110100110001110000000000011101000001010100010011000001000011110011110100110011111101110001110001110001010101010000001101001100010101110100111100000100000101110011111111110100110100001101000100010001001100000101110000010111011101000100110000011100000000111101,512'b00000000110000110011011111010111001100110101110000011101110001000001110100000001111111110000010000010000110101110100001100110001010001011101000000110000000000001101110101000100010000000101010011110000010011110001111100001100110100001111001101110100011100110001000101001101010111000000000000001101111111001101110001010000110001000011111100000001000000000111010001001111000001111100000101000101110101010100010001000001011111010011110100001100011111000111000111010100110100000111010111010001000100110000111111000111};
logic[2047:0]weight_l2[63:0]={2048'b11110000000101000001001111001111110000010000010100011100011111000001000000001111000000010000010011010000000101000011110000010111010111000100010000010001010011000001001101001111001100000000111101110000001111000000000001001100001101000011111111110111001101011101011101110100001100010000000000011111110001001100001100010100010000011101010011110001011100000101010101000101110101110001010100110000110011001100010100110000010000000101000001000111000100000100001101111111111100000001110000000101010101110001110001001100111111110001010001110101001111000000110001000011000011001100011100001100000111010100010111110000111101010011000011010011010000001111111100001100000100000000000011000011010011000000001101000100000100000000000000010100110000110000111100110000110001001111000100110111010000111101111111010001000100001101001101111101111100011111111111000101000011010001011111011100011111000100000000010001110011000000000000010000111100000011110000000011111100001111000111000100000001110101010101110100000001001100000001011111110001010101010111011100111111000100111101110000001100110000010000001101010011001100111100000000110100000011010100110011000000000001000000000011010011111101010101010001110111010100001100110001000000000000111101110101010000111101000001010011000000110001000101000011000011010101010000010101001101010111010111000100110000000001011101000000111111010000110001000001000100011101111100111100000011001101011111110000010000110011010000001100010001111100000001110011110000001111010100010001011101010100011111010100000001010101011100000011110000001101000101110000010011001111111101010111010011110011000101000000110100011100001100000111110011000011001111010100111100010000010101110000000001010011000001011100110001110001010100000011010001110011011111111101000100010001011101001111000000000011001100111100000011011111110011001111011111111100001100011111010100110100110000111101110001011111111100110101000100001101000000110111111100010111001111010001000011010001000101010001111100111101110100010100010100001111000001110100110101001111000101010111,2048'b01010000110001111100000001001111011101111111000100111100001100001100000001000000011111000001010000010111010011011101001101001111010001001101000100000100000001010000111100010001010111110001010000000000000111011100010000000001000111000000111100110011110101001111110000000000010000000100000000000011000011110100000000000101110011110011110011110111110100111100000001010000110001111101000001000011011100110000010000011101001101110000000001110101010011000000000101000011000111110000111100000011111101011101000101111100110100010000010111010111110001000101010101010111111101000000110001110011010100000001110000000100111111110111001100010000000001000100000000011111010100001111111100000000010100000100110011001111111111010001011101000001110100000101110111000000011101111100000100011100000001000011011101010000010111010000110011010101011100111111000101010001010001000100000011110111001101110100110001111101001101010011000011010000000011111101000111110001011100001111000001011111111101000101110100110101001100011111110101010001001101000000010111010001111100011111010011010111000111010011010101000101110011111101010001001101010000111100001101000101000111010001000001011111111100111101110011011111010111001100000011011100111101110011011100001100110011011101000001010001011101001100110001010000011111000001010100111101010011110101001111001111010001000001010101001100000001110100110001010001001100000011001111000001110000110011010001010011001100110001110111010101011100011101000001000011110101011100010001110001000011010011000101000000000101010101010100110001010000000100001111111111001111110101000101010101000001010001001100111100001100000011001111010101110101110100000011000001011101000100110001000100010001000000000001000001010001010001110111110001011111110011000011000011000100110000111101010100001101000001010000111101001111111101000101110011011100110001110101111111011101011111010000111111000001110101110000011101000111000011110011000001010011000001010001000011000100110001000111000011110000110000010111110011110100110100010011110000110011000100110100001101,2048'b00110101010000000011000000010100000011000001011100000111010101000111110000001101110111010001111100010001010011111100000011011111110001000000010000010101001100000101010000110111000100001100110111111111011100010100110100000101000001010000111100011101110001001100000101001111110011111101110100010100110001110111111100001101110011011100011101110011000000001100110000111111000011110100111100110001111111000001000111010000110101010111010101111101000000110100000100000111000100000000110000000000000100000111110111001111010011000100001111000011000111001111010001011101000011010111011101000100110100011100001100000100011101000100000111110101110000001111000011000001110001111111010001000000010000110111000101000000010011010111001101010100001100000111010111111111000100011100001100000011010001001111110000110001110001001100001100110101001101110101010001010100010101001111001100010101010000000100110000000100000100001100001101010111010000111111010100000111111101001101011111010101110000000100000000110101000000000011000000010001110011010100001101001111010001000000010100000001110001111111000000110100000100010001001111111100000011010101010001111101001111010100001100010100010100010101000100010101111100010111010111000000110000110000010000110101001100001101000101010111000101010100001111010000011111000111000101000101000101011101010100011101010111110000011111001111001101110101010001010101110011110011001101000101110001111100011100010011000101000101001111010111111101000001001101001100000011010100110100010000001101011100000000110111111111011100010000011111010100010111111100111101110111010101010011001100011101001101000011010011000101110111110000110011011111110001010001000011001100011100011100000111110011010011011111000011110111010000011111110000110011110111010000111100000111000101110111000001110111110001000000111100010011010000110101111100111100010111110000000101010101110111110100110111111101111100111100000000000000110000110111000111000111000100000011000111110011000000001100110100111100010001010100110100001100010101000011001100010000010100010111000001,2048'b00000100000000110111111101011101010101111100010101000100010011110101111100000111000101010100110000000000000011011111000000010011011101110011110011000101000000000000001100010001010000011111000001011111011101110000011111110001000101001100010000000000001111000100000011001101110011010101010000001111010100000011001111111100010001010101000000000101000000110000110100001100110011110100000011000111010000010100000011000101000111110111000101010100000001000101110000011101110100011101110011010000011100000111111100000011010101110000000101111100000100111100011100000111110001000111110000000011001101110000111100011101010001110000000100010011111101001111110011000000110000010111000011010000110111110000010000010100111100000100110011001101010100110100011101110100010011000000001100111101110101011101111100000111000000110111111100111111110100001100111100001111010000001100110011000000010011110111011100110001000001000101001111010100010011000101000001010011011111001111010011111100111100000000000000010000010100111111000011001111110111110000010111000000111100000001110101010001000001000001010101110011111111011100000100000100110100000111110000110101111100010101000101010000111100010011010000001111110000110101111100110101000111010101010000011101110111000101111111000000000100110101000101111101010111110011110001110011000111011111000101110100111101000011010000111111010100010011011100001111110100111111001100010101001101011101110011110011010000111100001100110111110101110011111100110000010101110100000000111101010011001111010000000111010101010000000101011111110101010011110011000101011101110111110001110000110111000001000001001101010101110111010100011111011111111101001101111101011111000011110101010101010001000111110100001101000001010001010000000001110000001100110101010100110111111100000100010111010101010000110011000111011100001111001101010011000100110011010100001111110001110100001111000011110011000100011100010000001100001100011101110101001101010100001100110011010100110000001101000000110100000011010011010100000100000000000011011100011111011111111111110101,2048'b01000100001100111100001111110101111111010100001100110011000111000100000100010100000000001101110101110001010000000000011101000111001111111101000101111101001111111101110101010011110111000001011101000100011101110011111100110111010101001100110000010101011100110111110100000111010100111111110111001101001111110111010000010011010011001111110011000111110100000111010101110101111100110011110100111101010111111111000111000011110001111100010111011111000101110011001111010011110100000101000000110101110000010011011111010101010000110001000001011100000000000101010000110100011111010000111101000100011111110111000101000111010001111101011111111111110111000111110001110111000100011111111101111100000100110011000000010001001101001100110001110011111100001111011100110100111100000000110000010101000011110000110000000001000001011101110111110101001101010011000011010100110000110000001100000001010011110100001101111111110100011101000111010101000100010000010101111111010001111111110011001100010001011101110011111101001111000011011111110111011101011101000011000001001101000101110111110000000000000011010011010011010000000011000000110000010100000011001100010001001100010111010100000011010000110011000001001101000111110000000011110100110000110000010001000000110101000100011100001111110000010000001111010100001101111111010000001101010001010001010001110101110111001101010101110000111100000001011111111101010001000101011100001100000000000101000101000100110011010001001100011101110101110011111101011111000101011100001100110111110001010000000001000000001111000100010100001101111101000001010101110100000011010011110111000000110001110001001101110101011100010000000111001101010011011100001101000101001111000001010100011100010001011111110101111111111101011100000000011100000000110101000000001100111101010100000011110011010011110000010000000001110111010111010111000111010100111101011101001111110101011101000100011100010001000011010011001111110101001101010101011100110101000111000100000111110101010100110000000000110100011100010100000001000101000111010101000001111111011111000111110101,2048'b00110101000011111100001111111111000011010000110001001111001111011100000111011100010011000011011100011100110000000001011100001111000000111111000001110000000100000100110011001101110111000000011111110000010100001100000100000000110001111101000101110001010000001100011100000001110011000111110001110111111101011101010111000001000101000111000000010101001100000000111111110011111111000001010101110000010011110100010101000100000001110000001100000001000011000100000100011111000101001100011111001111010011010001110001010100000111011100111111110100110011000011010011010000110011010011110011010101110000000101010001010001011111010101010001111111110100110011110011010000110000001111110111111111110011010100010100000001110011000011110011110100010100010001110101011111000000000100110111111100110001000101110111000011000000001101000011000111000001011101011111001100000100001111111101111111001111011101010000110000110101010111010001110101010011110100110011110001001101110101111111010011001101011101001101000101111101000100011111110000000011010011000001001111000100010001001111000100010101000101000100111100001101110000111101111100111101110101011101011101110111111100000001110000111100111111010111000000000101111101110101110100110000011111000101010000001101111111001101110111110001001111110100010000010011010101110000000000000111111111111111001101010001110011000011110000010100110111110101000100011101010000010000000011110001010001111101010000010000011101010101010001000001000001010000010011011111000001000111000101011101011101000001000100001101000111010111000000010000000011111111110101010101010101111100000011110000000111000101000000000001110000111111110001010111110001111101000001000101000011011101111111011100001101000000110011111111110001000101000011110111111100000011111100001111000001000000110101011111011101010000111111010001010100111101000011001100010001000101001111110001010000001101010111111101001101111100110100000111010101010000110011000000000111110000011100110001001111000100001101001100110101000011000111001111110001110100110100010011001101000101001111,2048'b11111100001111010101011100110000011101110101000000000011111101000001000111000000111101000111111111110000110100000000010001111111001100011101010000000101110101010011111111000111110001000001000011010100000111010011110000001101001111010001110111010011110011010001010101111100110100111101000111010101010100111100010111000100111101110000010100000111010000011100010000000000010101110011110000011100000100111111010001110111110011011100010011000000000111111101001101110111010011110000010011010100110011000100111100011111000011010011010011000011110011111100010100000001011101000111000000000101111100000001111101111100000000010001001101110011001111110111001100011111010001000100010011000100000100110000000011000001011100011111111100110001001101000000000000110100001100110100000000111100000100110111011100000111000111011101011101010101000100010000000001110001011111001101110001001101000100000111110000010100010000010111110011110111000011111101000100110001000000010100001100001100000101010001000000010000111101001100001100000101000011000111010100010000000100110001110000010000010100000011001101110000110111011100011111010000010000000000001101111101110100110111111100000011010000011111110101110111000101000111000101000100000000110000110001000001110000110111000011010111110001000111111111111111011100111100011100010111110100001111010100000111011111000001110000010011000111110001000001001101000111011111000001010000011100010101110011000011111111011101001100001100110000010100000100000000110101110000110111000111011101000011000000011100110011000001000011000001110011010000000100010111000000000000111100011111111101010100010001011100110011011100010100010001010000000000011101001111000111000100010101010011000011000011110011011101001111000100001111111100000011010101010100110000110011010011010101110101011111011101111100110011000011111100011101001100110011001101000101011100110001110001011100000101000001000101110001001111010100111100010001110011000000011100000011000001000011110001011101111100010111000100000100001100010101000001010111010000110111110111000011010001,2048'b01010000010000110111001100011111110011010111110001001111000001000000110000111101111111000111010111000100000100111111000101010111010000010100111101110001110000001111000111000101110011110000110000110011010000001111011101001100110111111100110011010100001100010011010111010011110100010011000001110101110100110000011111010100111111110100011111110001000001011111010001110000000111010000011100111101000100000000010000000111010100011100110101000100001101110111110011010001001101001100011111001101000101010011010000110011010000000011011101010111111111010111111101110111000001000000110111111111110001001100110000000101000100110011011111000100000101001100110111000101010011010001000000011111010000011100000000000000011100110111000000010101001101001100110100001100000100111101011101010001000001110001000100110001011101000111111100000101010100000011110101010111000000000001110100001101000011010000000001000111111111010111010001000011001100001111000000111111010000000111000100110101010000000001010011000001111111000100010000011101000111111100000011010000000111001100000000110101010011111101000011000101010011011111010001000011110001000011110001001111111101000111011101111101110001011101000000010001000011111111111100010000010000000001000011000000001101110111110101010011110011000000010011001101000001000111011100110011001100010011010101110011001100110011110000010001110111111111110101010011000000110100111111111101111111010001010100001100001111001101111100000011001111111101001101000000010001000111001101010000011101110111010011110011011101110100110111000011001100000100110011111111001111110100110001011100010011000100010101011101000011110011110111010111110100000100000000110000000001111100010000000101110000111100010011010011010100000111110000111101010011011100001100110111000000000101000001000011110111011101111100010011110100010101011100001100000001110001110000010001011111000011110011001101010011110000110111000001110111001100001101000000110000000111110111010101011101000011010001011101110001111100110000010100000001000100000100010100000111110100001100010100,2048'b00110100000000010000010101010000110000000111000000110101010011001111011100011111001101010001110111011101011100010100001100110101000001110101001100111100011100000011000001011101110100010011011111010000010011010001110100110100011100111111000111000111000101001100110111001100001111001111110111110100111101110000110000110100000101001111010100001111000000001101000001111101000100010111111100000111010011001111000100110111010100111111010101010100110000110000010100000111111101000100011101010101111101000000000100111101000011010101110001011100000000110011000001111101000111110011000000001111110111000011110100000000010001111111000011010100110001111100110100000100110001010101010100000000110101000000000100001100111101000111111111001100000011001101110111010000000001110100000111010011010101010101110111000011000011111101000011011101010001010001001100110001000011111111110101000111110011011101001100010001111100010101010001010100010011000111110011110000000000010100001101001111111111001111001101110001000000110011110101001100001101010001010011010011111111011111011111001101010101110111000100010001110000000111111100110101000100011101111101011111001100001101001101011100011100110001000111111101011111000100010111110111010111001101000001000001001100000001000011010001001100000000111100010101001100011100110111000111000000010101000000000001110100011111010001010101011100110011111101000001010001011101010000111100000100011111001100000001110100110100010100011100000111000000001101110000110101111101001101000111000011000100110011000100010111000011110000010001000001000001000111111101010101000011010100010100000000110001000011000001110000000001010111110000000100011101110100111111110001111100010011000101001101111111000000000000000100111100110000000100110100001100111101000101000000010011010000110001000001000100010111011101001101111101000100010001001111110111001100110101001100111100110111001111011100000001010011110100110001010000001101010000110011011100000000110001000000000100000001010001010000000001001101010011000000110001010101001100010000000100110001000011,2048'b00110111111101110000110100001100111101011100000000000000110001000011010000010011110100001101000001110111000011110101110000110011000011011100011111010111000001010100111100110000111101010000000100010001010100001111010001001101000000000101110101000001010001010100000111010101000111110001110101110001001101000000111100010001000101001100111100000011010000000001000001000111010000010111000000111100000001011100000111010000000011010011011101000001000111110100111111000100011101010011000001111101110000001100110111000011000111000011110001110100000111010101010000110011010101110100010111010111000111011100010001110111110100110111000111000001111100110101010111110111010001110011011111000111110111110011110000001100000000110001010111110011111111011101110000010001010001000000011100010100000101110000110001001100010000110101011101010101011101110001110101010111111100000001110001110001000100000111001111000111000001011101010101001100010011110101010111110000110011001111001100000100110011010101000100010100110001010100000111000000010011001111010011110001001111010100011100011100111100010100010101110100010111110011010001010000001100110001001101010001110000000000110011010100110011010100110111110101001100011100000101000000000100011100010111000011010101111101010000001100111101000000000000001100001100010111110111000000110011111101110001110101111100010100000000000000110101010101001100010000000000001101000000011111110101000100110000011100000001000001011101000100110100111111110001010100010001110001000100000111010011000101000100001101000001010001000101110011000101011100000100110101001100010111010111010000010101111101110111111100010101011101010000000100011100001100001101010111000011011111000100000101000111010100000000000101010111110000110101010100010101000111000011011111000001000101000111010111000001000011001101011100111100000011000100010011010000001111000111010000011111000000000100000111011111010111010100110101111101011101001101110101010100000000110001110101110011110111110111010011011100010111110000001111001101000000011101011100000011000100001111001101,2048'b11000100001101110000011111110000000000011101111101000111010000010000010001010001001111000011010001010011111101110100000000000000110101111101011101010101111111010001010011010001000100010001110101000111010001001101000000011111000111010001110011111111010101000101110111000111010001010000110101000001011100011101011101010001010111110111110001110101110001010101110111110100011101110100011111111100110001001111110011010001110101110001010011010101110001001101110100111100010100010000011111011100001111111111001100110100011100111100110000011111010100000100111101111101000100011101011111111111000100010011011111110101000001001111011111110101110011010100001100001111010001110000110111010101110000110000000001000001110011010001000111010100010111000000110011110101010000000000110111000100110000000001001111000100001100010111110000000000011100010011010011001100010111000100000011011101000111110100001101000000010011011100111101111101110100111111110101110001011100111111000011010001010011110100110001000100000101000100011101000011110101010000010001000001001100010101010000001101000000001100000111010111110101111101111100000000010001011100000100000011000001000111011111010100010111000001110001011111010111011111000000110101110011010101110000011111000111011100001100010111001100110000000111010000011100000001111101110001110000110101110001000000010011000000110000001111110000110001111111000011110100111101110001000100111100000000000100110100010000111100001100010101010101111100000000110000001101110011110101011101011101000011010100000111000000000000010101000111011111000001010100010000010001001101010111110100000111000100010011000011000000010000010000000101110011010011011100010001010001011111011100000000010000011101000001010101011100110011010101000000011111011100110111000101111111000001110100001111010000111111111111011100010111001100110100011101010000110101010100110000011100000100011111000111000001000111010011110101000011011100000011010000010101010100110000010101111111010111001101110111011111011111000100000100000001000101110001000001001111011111000000110000,2048'b01000011111100011111000000110101001101011101010000000000110000011100110011110011011101110000001100000011001101111100111101000011011100010001111100001100010100010011010000000000010000000000000111000001010000010101010111001100000000110011010101110000110011010101111100110100001111001111000100000100001100000111010000110011000111001111000111010001000001000101110000001111110101110000001100000111110011000011000111110111000111110111110100111101000111000100010101000100011100111100001111110001010111001111011100011100011100110111001101001100010001110000110100010100001101110001110000001111111111110000011101010100000001010100000001110000110101000011110100110011010001000000001101011111110100001100010100011100001100010001000000110100001111000011000111010000001100010001011111011100000101110100111100110111000011011111000101011111110001000011001100000011010001010100000111000011000011000000110001111101110011001100011100011101000111010111111101110111010101010111000100000000000000010001000001010000010000000011011100111101011111010000000100001101110001110111010101000011011111010101000001000101110000010011011100001101110000001101010001000011110000111100110101010011010100110000000001110100000000000111011111000101110100010100010011010011000000011101000100000011110101000011000000001101010101010111010000010100000111000011000000001100000001001111111101110100000100011100111100111111000001111101001100010101011111010001110100111101110000111101000011000001011111110001110000010000010101000101111101110100001111011111111101010011110001001100010111010011000100011100000001111100001100000011010011110000000100001111111101011100011101010000000000000100010011110100001100001111001101001111111101110111000001000111000100010111110001110011010000010101000101000011010011111101110101010000110000011100010001000000010111010000000000000011000000000000000111000101011101000011110000000100110011110111010000011100011100011111000101110101000000000111000100010011001101000001010100001100001100110100000101010001010111110101111100110000010101010001010111001111110011110011,2048'b00111100110000010011011111011111001101011100000001000111110011110101010000110011111111011100000111000011000011110000010000110100011101001100010011000011011101000011110001010011010100001100110101000011001111110001111111000011110000000100001101010111000100001100110100110001010011000000000100010000000000010000000000110100010100000100111100001111110100011111001111000100010101011100000000111101001111110000011100000000011101111101000100110001110100010101001111000001010100111100000011000000111100011111010001001101010100000000000011110001111100110000000000010000011111000011011101110101111100011111000011000101001111010111111100111111111111110000010000110111010011111100010000110000000011111111010001110111001111010011010011111100010101000101010100000000111100010101010111010111000011011101000101000100000001001111000001011100011100110100000001010000000101000001000011000111010011000001110111110001111101011101010101000000001111110000001100011101010100001101111111010011000011000011110011000111000011001100111111000111111100110111010001110101110100000111010100001100110001110011110001111100010001110111001100010011111101110011001100000001000001000011110101111111000101000001000011011111010100011100110001000001000100001100010000001100111100000011011111010001111111001100011111001100110100111111000001110011011111011100111100010000110000001101110111110111010000010001010101001101000000000111010011000100110011000000000000001101011100000100110101111101010000111111011111110111110101001111111100000101011100010001011101001100011100010111111111111100010111011101000111000001110101001101010011000011000000000000110100111100111101001111010001001111110011010000001111110101000001010011011100000001010001110111011100010000011100110111010100011101000000110011000000001100110100010011000000111100010100011100000000000100000011110000011100010000010001110100000100010001011111001111000001001100110101111100001111111111000000010011000101001101000100011100000000011111000000111101010101110100111111010000010101010001011100110111110000000011000101000100001101110000,2048'b11111100110000000100010001011100110101110101000111000001110100111111110000000001011101011111111100011101111100000111110100010111000001011101000000000001000011110000110001000011000100110000000001111100110000110101111101000111110100010000000001000111010111001111111100000000110000110100111101000100111111110100011100110111110111001101000001010111010111000001110101000111000100110000010101110100010001000000000000000011010001010100000000000000001100110101000101000111000011111111011111010001000000000100001101000101111101001100110111000011010001110101000000011100110101011100110011111100110001111100000011111100000111000001010000000001000111110100011101010100111100011100000101110101110000000001000100000000110111111100011111000111110100110111011100000100110000001111001101000100111111011101011111001100010011001111000001000101000001110101110000000000111101000100011100000001000111110011000000000000000011000011110001010000111101110111110111010000000101000000010000010000110001000001000100000011110000011100110001000001110011010011010111110000110001000000010111010011000000001100001111110001110100010001000000011100010000011101111111011100110011110001000111000000001101010111011100111111110000000100110100111100110100010100111101000000010001001100110101011100010000010100110100010001110101011111010000001101001111001111011111010101010011010100000001000011010000000100000100001100001100010111000000001100000111110001000101010000000000000111110111111111000111010101011111001100010011110000000001010111111111011101010100000101000001110000111111000100110000110101011111110001010001000111001101000100010011001101010000110101110101111100111111010011001111010000011101111101111100010111001101000011110100000001110001110101110000010011111111001101000100010000000011000111000001000000001101000001000111010000010100110001111101011100010111010100000111010111111101110000001111000000000100011101000000010100110000011100110000001111000111110000010000010001000011010011010101000101000100011101001100000011110011111101111100001100111111111111111111010100110001010101,2048'b00010000011111010100000100001111110001000101000001000000011101110001110001110011110011110001110011110001011111011111010101010001110000010000110011000011110000000111000001111111000000001111110000111111110100000000011100000011110100110100111101010011110000110101001111111100010101010100011111011100110011111111000011010011001111000100000001001101010011010001000011110001111100001111110000010001110101010001000101010011001100011101010001110101111100010011010100000001000011000111111111011100010001000000111100110000010000110101000001010100010011111100110101000001110000001101001111110011010111010101110000000101000101110011011111110111010111000111010001111111011100010000010100110111001101111101110111000000010101110001011101110000010000110001111101011101111100111111010000010100010000001100000111011101010001000011110100111101110001000011110101000001000100010000110100010000001111110001000000000011011101000000110000000111011101000000001111010111010011010001111100000001000001110111110011001100111100010000001101010011010000000000110100000011000011110100110000000000011101011100000000111111110000110011010100001101111100010011110101110101011100011101110000011101111111001111000100010000000011010111000100110000110000111111001100000011010000010100000000110101001100010111010011110000111100110111000101000111110000010011000111001100111100011111110001010011011101110011010101010001000000000011011111001100000100010001000000011111111111000000000100011111010101000100000001000101000100010100000111001100010011110000000111010011110000000111110000110011110111011100010100110111000101000000000001001101011101000011011111001101111111001101011100000001001100010101010101110100110111001111111100010101001100010111110011000011001100011100000100000000010011110001010011010011010011011111000101011111000011110001011111000100111101000111001100110011110100110100001111010000000000111111011111110100000111001111000001001100000001000101011100010100000100010011000011110101110101011100010001000000000001000111110101001101000001010100110000001111010101001111001101010000,2048'b11010111001100010011010000011111110011110000000101110000011101110101111111110100010111010111000011110011111100111100010100010001000001000000110111000100110111011111001101110101011101110100011101011100000100010111010001001101010101000001010111010000000001000101010001110000010000001100000111111100001101000111110111110101011100110100111101000011000100010011010100000100010011000000001101110101110000110001110001000011001111001111110011110101110011001111011100010101010101110000000000001101111100000011001111110111110100000001110111111111010001011111110100110100001111110001011101001100000101000000001100110000010100110000001101000011001100001101110000000101110000001100111101010111000011010101011111111111110011110100010001110101000000000101010011000101010001111111111111011100111101000011110001110000010100011111000101110000110111000011110011010011000011000100000011110001110000111100000011011100010101000101000100011101110000011101010001011100110111111101111111001111000000010100000000010100010001011111111100011111000101000111000100111101110001111100000001000111001100110000111100011100011101010001000111000101110000111111000101010100011100010000000101011101001111110111010000000000010001010000010101001101000001110100000000011101000011000101010000011101000000110001000011111111000111000001000111000011010101010101111100111101110111010111001111010101001111110111110011010001010000010001000011110011110000010001110011110001110000110100110011010001010011111101010011010011010101110101001101110000000000110111000111010100111101000000110000000100110000010101010000110100010001000000000001010011010000000101000100011101000111110000111111000000110000010011000101010011110000001111000011011101110000000000011101010000110100010000001101001101000000011100001101001100010011000100010011011111000011110111001101111111001101000111010011001111000000010001000100000001110000011101000000000000010111110101010000001100110000000100110000001100110101010001000001110011011111010101110011110011010001110001011101010000111101110001000111110011000000010101010011110011,2048'b01000011000111000100111100111101011100001111000111110011010111000001000101110000111101000001000111110000110011110111010000110111110111010000010011010000110111000011000111110011010111010000001111110011001100011101000100111111110101110111011100000101110101000101010111110111001101001101011101110000010101110111000111110101001101000000000100000101110101110101001101110001111101110000110000001101110011001111110111001100011100110011001100000000000100001111110000000011010000110000001111001111000111010100010101011101010111110100010000000001000011000011110011001101110000000000110100001101110000001100010100010100110001010111000100000011110111000011000011000100110001000011110100011101010000011101010111011111110101110101010100110011000011000001000001011111001111000111011111010101000000001111001111000111110001000000001100011111001100010111111101000011110100011101010001000000000000001100111101111100111111110000011111011101010101111111010111011111000001010101000100001111000100110011000111011101010111111111010101001101010100111111010000000001010011000001001101000100000111010001110011010101000101000111000100000101111100110100000011000101110011110001001101011111110001011100110000011101011100110000111100110011110111111101010001010101001101000000110001010001010011000111111111010111001101111111011101111101000100110001000000001111111101000100001100011100001101111111001101000001110100000111000001110101001100000111000001000011011111010000111101011101110001000000010000000100110001011100000111001100010000000101001100011101110101000000111100000011000011111111110111010100010000000100110011001111000000001100010111001100011111010011010111000101011100000001111101001100000000011100000100000100000100010000111100110101010000111111001101111111001101010000001100000111010100110001011111010111111111000001110111111111001100010100111100000000001101011100000100111101011100011101010011010111110000001100010011110001000000000000111101000001001111001100000011011101000001010011110100111100110000111101110011000000000100000111000001000011001100000001010000110011,2048'b01000000001101110000010100000011110111110000010100110000111100110011000011000000010100001101000001001111110111110000010101000100110000111101110100000101010000110011000000110100110100000101010100010000000101001100011101001111000101111111001111010101011100000100000011011100010011111100000000110111110011011101110100000011000000010100000111000100110101000011000111000101010000110101010000111111010000000100110000000101010101011100000011010001010101010011000100010000001111011101011111110001000100110000110111000100010100010001110111011100010100000011110101000100110011000001001100001111110011011100011111010111110001000000000011010101011111000101000011000001000011010011010101111111000100110000000111110011000111110100000011110011000000000101110101010111110111010000011101111100110000110000111100011100111111010000000100001101001100010001000001111100011111110011000001010000001100110000110111010111001100001111000100001111010111000101001100110000110001110011000101000101000011000100110111000000011100010100110011110101001100110000110111001100000100001101000011010011110111110101011101000000000000011111110100010101000011000001110001010111110011110000000001001101010111110011010001000001010000001100110000011100010111011101111111001100110101001111000111010011001111001111110001011100001111110000111111001111111100010100111100001101111101000011110011010011110101010000110000000000011101001111000101001100110101001100110111010001010100010000000111010111110001000000001100110000110001001111000111001111000011000011010101111111011111110000110001110001000011111100001101111100000011011101001111000001000111010000011111110111000101001101110100000111010100110111010011000111000011011111110100011101001111001111111100000001010011000111011101011101110000111100010011111101110101000000110100011101110011010001010001000000000000110001111111110011001100001100010000000000111101110001110001110011011111000111010011010000010100110100000011010001000000011111000000010001111111010101011101110100011111110111110100110100001111000100011111001101000111111101110011000011,2048'b01000011111111110000000111001100110100000000000001011100010000000100110011011111000000010001110000010011110101001111000101010111111101010001110111010000111101110111010100010001010001010101000101000111111101000001110011010100011100000001001101010000010001111111010000010000010001010000111111001100011101010111011100000111010101110001011100110000110001000111011101001111010011110011110101010011010001110011000100110011110101110111010011111100010000000011110101110101010101010100010011010100001111110111000101010101010000110011110100111111011101010100111101110000010100110011010001010011111111000111110001010101010111011101011101110111010111000000110111110000110001010111000000010111111100010100011101000100000000110011001101011100010001111100010000110101000011110001011111000001000001110101111111000011110011000000000101000000111100000000000011111100000001000111010100110101011100001100000000001100010000111100001101000100000000010000011100010000000001110100000000000101011100010111110101001101111101000100110011000101010100000011010101011111010111010101010100010001011111110111000100011111000011010100001101010100010001111100010100011100111101010101111100111100000101111111010101010000110001110000110101001111011111110011010011110011110101011100001100011111010100110100111100011111110000001101001111111100000011110001001100110100111111010011001101010000001111010111110111000101110100010011110000000000110011001111111101011101000000001101000001010011001101110100110001011111110011000000110111010101001111000000000000000111111100110000001101000000000100000111010011010011000011010101001100010101110011000101000111000100011111110000000100110111111111110100111111010001110000111111000101010001000000110000010101110000110011000011110100010100000111011101000000000100111111000011001101000001000111000001000100110100000001000011110100000011010100000001010000111100000001111101001100010011110111000011001100001101000000011111111111010000000100010101010011010100010011011101111111010000011101000000010100010100110100010000110000011100110011010101010101010100,2048'b01110011010001110101110001010111000101010000111100001100000111011100010000110001000111110100011100010001000100010100000100110011000001011100011100010011110101110101000000111101000011110000001101110011000000110011010000011100010100001101010001110000001100110000000011000111000100000000111111010101000001011100111111010100010100000101010000010100110011001111000100000100001100011111111111001101010000000011000011001100010111000011000001000000110100001111011100110000010100111101111101001100111111001100000100010100000100000100010000011111011101110011110000110000001100000011000011011100110100011101000111000001010100111111000011010101011101010011111111001101001101010011011111000101000001000001010111110100000000000000110100001100110001011100000001011101010011000111000001000101001100010100000011010000010111000111001100010001000100110001000100110011010101110101010111000011010111011101000011001100010111000001110100010101000100111101000101010111110001110011000011001100000000001101000100010111000101000100110011011111000111011100110011000011010001000111011100001100000001001111110111110101110111011101110000011101000101001100000111111101000000110000111100111100111100000001110100010001111111111111000001010100110001110100111111111101111100111100000011001100001101111111010100001100000001110100000000110100010001001101011111010011010100000101000100000001110100110111001111000000010111111111001100010101000000111111010000000100001100110000000101110000010111110111110011010100000111111100010000001111000111110001010000001101000101000101000100110011010101010011000000011111110001010111011101000000110011001101000111000000000100000001011101001111001111110111011111010100110100011100000111001111000101001101001111000111010011010101110000010100000011000000000100000011110011010001110000111100000011001111110001010111001101010100000001000011000111000000010101110011001100001111000000000011110000010111000101000001110000010101111101001100111111000001110011000011011111001100011111110011110111000011110001011111011101111100000101000001110101000101000001010100,2048'b01001111010000010011001101111100000000010011110000010011110001111100111101000001001111111100111111001100111101011100010001010100011111111101110101110100010000001100001100110100000000011111110100111101011100001100000000001101010000110101000100011100111100110011010000010011000100010001001100110011010100001111110000010001110001011111000001000011110000001111110101010111010100000000000001010001000000110000011101110001001111000111000101000001110111000001110100110101001111010001110100001101010100110100011101010011000011111100010101111101001100110001000001110001000000010001110111011101111100110011000101111101001111110101001100001111001111000011010100011100010101110011001101010111110101110101001100000111110111000001000011111101110001000101000100111101000001111111000000010101110001001111000011001111111111010111110001110101010101110101000100000000010001000100111111011111000111010100110000000100000100000100000100000111000111001101000000111100110011010000110000110111110100110001111101110101000000000101010001110011111101001100010001111100010011110000110001010000110011000000011101011100011111110001011100110101010101110100110000011111110101110100011111010100010101010101000111000101111111000001000001010111010111110001001100111111010001001100110000000101000111010011000000110100111101001101000001001101010101011100010000010111010001010100001100001111001111011100110111110100011111010000010100001100110101000000010011000011001111110011111111110011001100001100011101011100001111000101111101011111001111110100000001000001001100001101110000001111110001110000110011010001010000001101010100000011111111010101000000110000010000110001011111110011010100111100110011000000110000110001110000000000010001111100000011000001001111000111000001000000010100010011001100110100000101000001010000110011010000111111000011000001000000110100011101010001010000111100110111000100001100110100000100001100110001010011000000001101000100111100010011111111010111110001010101000101010000000001010001000101000011001100010100110101010100000000111100110111110001000001110100000100,2048'b00010111001111110011011101000011010001001100010000110111000011000011001111000101000011111101000101010001000101000011110100000101000011110001000101111100000101001101001101000011111101000011010000001111001101110000001111001100000000000111010101110111011100011101111101110100111100000001000001110001010001000000110011110100110100010011111111001100110011110000011101110100011101000001111101000101111100001101111111000001110100000100000001000011011101000100000000110001110011111101000011011100000000000001001101110011000111000101000000111100110100000011010100001111011100010100110001000001110100001100001111110000001100111101001100010000111100000000010101000000011100010000110001111101010000010001000100110001001101000100111101010000001101011111111100010111010001110100111111010100110111011100110011001101010001001101000001010100011100001111010001000111110100010001001100000101000101001101110101010000000101001101010101110100000000010100110111010000000011000011010000000111110111111100110011110111011101010011000011110000000000110111010111000100010011110000010101010001010011010001010100000011000111011101000101111111110101000101000001011101001100011101000100001100110100110111010100001111110000010001000100110001110100011101011111110101111111010000111101010011111100110100110111111100010001010100001111000100110001000000011100000100000000010101110101000000001101001100000111111100010011010001001101010100000000001101011101000001000100010000000101010001110011110001111111111111110011001100000100010011110001110001010100111111011101001100010111110000110101000100110101001100110000010001010111010011010101000011110001110011110000000101001100001101110001010000001101000100110100000011000000010000001111001101000100110101110111010000010000110111000001110011001100000100110100010001000101001111000011000000111111010100111101000101111101001100001101001100110001010100011100001100001101001101000111011100000111111101010001110101010001001101011100110111111111011101001111110001011101000011000001010111000001110100001101010100011100000101111100011111010001111100,2048'b00110011111100000100000101010001010001000100010000001111010000010001000011110011110001000000000100010111011100000011001101111101110000010011011111000011001111010100010111000101000100010111010000001100000011001100001101000111110001000111000101111111000111000000010111000100111100111101000000001100001100010100110101111101010011001100000001111101111101001100111100001111111100010011010011010011010000000000110011011100110101010000010100111101010000110100000101000001010001010011010000011100110011010111001100000100110011110111011101010100010011010101110100000111010101111111000000001101011100010111110101000011110100000000000100001111000100110101000100001111001101011100111111010111001100000001110011010000011100001111010011010000111100000011000101001101110100001100110011010011000011110000011101111100000011001100110000111101010011011100110100000001110011000100110011000101110000010001010011010000111100000111110111111111110101010000010011110000011100011111110000000000010000001101011101010000000111000001000011001111000001010100111111000001110011011111001100001100011100111100110100001100000011000101011111010000010100000100000111000001011101010101110000110111000000000101110101010011000101001101010000110100111111001101001111011111000001110000110011010100000111000100001111000011110100000100010101111111000101111111000111010000001100000101000011001100000100010011000100110011000111010011111100011100111111111100010011011100000011001111010100000111011100110000001101010001010101001111110000000011000100011100010100010000001100000100011111001101000001110111010100001101111100010000001111000101010011110111000111111111000001011111010001111111111100001101110000110101000001011100000011010101010001111100000111010111000000001100000000010000001100011111010001010011010111110011010000011111010111111100001101111100001100000111000111000100110100010001000100110101110000011111011101001101010111001100000011110111001100001111010000000000011100010000000111000011000011111100110011010100111100010101000111110100001111110000111101110100010000111111010100000011,2048'b01110000111101000000010001000011010111110101010000000000110011110011111100001111001111000101000101010011000100000100000000010000111101010011001100000011000011010100011111000111000011010011000111110101010011110111000000111100111100110001110101110011010001110001110000000011011111000001000001000011011100000100000000110000010001111101010101011101000001110000010000000001000100011111010000001101010000001101111101000001000011010011000001110001010101011100001101000011000000001100000011010000000000111100110001000111010000010011010001000001111101011100000100011101110101010011011100111101111100110100011111010011011111110001110000000101110000111111000111111100110001111100110011001101110100011100001111110100000100010100111100001111000011000011110101000011000111110001000111011101010101010100000000111100000111010001000000010000111111110111011101001101110000001111110001110101110011000011111111110000001101110000000000010101001111010100001100011111010101010111001111111111000111010100000111010111110000001100011100010011000111000000010100110111010011111100110000000101000011110101000001010001011111000101110101000100010001001100010000110111010100000001000101000111010011111111000101000000111111010101110111010000111101111111000011111101000101001100000101010000001100011101010011000000111100000111000011011101010100111100110011110000010111010000010101000000010111110101001100011101010000110111000101110011000000000001000100011101010111000111010011110100000101110011011101000000000001110011011101010001110101110100110001010011010000110111001101000011110100000111001101010000110011010011111101011111000001110100010011000101011111010011110001111100011111111100110000000001111111010101010000000011011101001101001101010111001101110011000111110100110000110000000100010000110111000011011100010001010000111100110001010100000011001100000001000011010011000101000001110101111111010000110011001111111101110011110011000011110001110011010001000001011100010000010111000111011101011111110001110001110111010111010100001101110100110011001101110000111100000011001111001111,2048'b00000101111100111100000101110001001101011100010000000111010101011100000101000011000011000011001111111100011111000011000111110100110000000111011100110000011100001100110100111111011100001101010100000011000001000100001111001101000111110011001100010111010011011111000000111101111100111111010101010101001101001100110111110001111111000001010000000000000111110101111101001101111101001101010100110001010000010000110000110101010000000100001101010101000100000101011100110000111111110111110001001100110000010000010100110111000000001111010011110011001101001100001111000100000001000100110011000101011101011101110111010001001111110111000100000101111100000011000000000111001100010001010001000111001111000000110111011100010011000100110101111111010001111101111101010000001101000001000011110000000101011101010011010000000011000011001101110001010011000000111101011101111100111111011100111111111101010001110011001100011100011111011111011101010111010001111100000100000011011111110011001101010000000000010000000001010001010011001111110011110000010101010011111111010001111111000001000111110001001101000100000001000100111111000011110011000011010100110011110101000111110011000000010101011100110000011100010000010011001101010000111100010011001101011100011101010000000000000101000000001111011100000001010111010000010000011100000101111100111111001100011111010001000000000111000011010111111101000100001100001100111100111101001101110100110011110100000000000100000001010001111101010101001100000000111101111100001101110101110001110011000000001101011111110101011101000000001100000001111100010001110001000111111100001101110000011100001111110000000000010101010101111111010000001111010101110101010000000001110011000100001111000100110111111111000101110001000100110011111100110100110101110100001101110101000001000101110100111100001100001111001111111101010101011100001100011111011111010100011100011101000101011111011101110100011111010000011100010111000111001101110001011101011101010000000100110111001101010001110000000101001111011111110001110100111101010001111100011100011100000011000111,2048'b11110100000101001111000101010111011111010100000101000000111111110101010100000000001101111100010100011101110000110000001111110000000000010011000000111100110111000001000000111101000100010111000001000000000100011111110000111111000101000001000000001111110000000000011111010011110111110011000011000000000100010101000101110101111100111100010111010111010100110100110001111111001111110011001101011100111111110011110011000000010111110000110111011101110001011111001101110111000000110000011100111101111101110101010011010100001100000011110001010001010101011100000001110011000000001101011111010100000100010111010001110100000101111101000011000111010101111101110111000111110001001100010100001111000011110000000000000000011111110001000000010000000100011100011100001100011111010100011101000111111101001101010100010000110111010000110100001101001100110000011101000101011101000100001100110011001100110000111111011111011100000111110111010000001100001100010100001111010111001100110000110011111100000000000100011101110001110001000111110100111101010001001101000100010111001111011111110001000011110011000101000011011101010000000111011100110000001100000001000100111100011100000000110101111111001100000000000000011111001111000001001111001111010100110000000100000011001100000101010001000000000011011100000011000011001100000001001111010000000001001101001111010111110001011111010011010100000100010111000101010101000100110000011100001100110100011101000000110001110100011100110101011111110101111101110000000100110000111101001100110001001100000100111111001101011101011100000111001100000011001101010000000011110111000100001111000100000101110000010100011111010000111111001101001111110001001111010001000001110100001101111101011100010100011111010001111101011100000000010011000001000000010000010000000100000011000000001111011100110111010100111101001100001101010000110100110111111101000111000100001100001100111101010011010011010111110001011100001100000001010101010000001111000101111111110111001100110111110100000100110001011111011100010000000000000100010000110100110000110101010100110001,2048'b00010101010011000111001101110111010100000111010111010100001100011111011111000111001111110111111101010101010011000011001100010111010011010001110100111101011111011100011111110111011100111101000000000101000000001101001111001100111111001101011111000101010101010101001100010001110011001101000101010000110001111111111100000001011100001100011101000011010001011101000100000001001100000011010000110000010011000111000101011111000000010111010101110111000111001100110000010001010000001100110111011101010100000011000000011111000100110011010100000001110111110011000101010111111111011111010000000100000100011100110001001101110011001101011101000000110000011101110011000011000100001100011100110011000101110011111111010101111100000101000111110000010001010111110000010100010011010101000100110101011101010101000000000001000001110001110111011111010001110001000001110111000000011101001111110100000101110001010011001101001101110000000011001101000000110111001101000001000111001101010001010000010011010000110101001101011101011100000000110100011101110111010001111111110000010101010001000100111100111111010000110101010001000011000111011100000101011100001101000011000000110011001111010011111101110001001100111111011100000011010011010101000100000111001101010000110001001111011100010000011111010000000001000100000011011101110111110011010001010011110000111111000000110100110000110101001100110100011101010001110100110011001100010100110000000001111100110011001100110000111101010000000000011111010000010011000111110011010001110000010100000111010100011111010001110000110001011100011111010111010111010011010001000011000101001100110011001101010000000000001111001111010111010101001101000011010001000000000100010001000011010011000011001100011101001100000111010101001111000011011111001101010111110011111111000001010000000011010011110100000000000000110100010000110101000101110011000111000100011100000001000111010100110111010011010001110000000011110101011111010111011111011111010111110011001100110000000011000011000100000111001100110001110111111100011111010000010111010011110001001101110101,2048'b00000100010111000100010001110111000001011100010001001101011101010000010101000011110111110000000000111100000001001101110000001100001100011111001100110111110001001101000101110011010011010011110100001100110011011111110100001100001111110111000000010011001101000001000111000000001100000001000000110100111101000100000011010101001111011101000000001101111100110000000000110011000111001101000001001100110000110001111101111100000100000100111100000101000111010000000101110001011101110011000100000000001100011100000001000000010011001111001100010100011101010011001100110011000000011101001100010011110001000011110000011100001100110000110011010111110111011111011101110001010011000000001101011111111101110011011111000000110000011111000001110111110001011111110101110000111100111101110011000101110001111101110100110001010011111101110100110000111100001100000001000000110100010000110111000011000011000000010000000011111111110100001100001111010101111111001100010001111101011100001101110000010001110000001101110001010011000000010111010001001100110011011101110100011100010100000111000011010100110000111101111111010001111101001100111101011101110101001111011111110100000001010111000101110101110001011101110100011111011100010011010111011100110111011101001101111101011100011111110000110000110100111111010000000101010011010000011100011111011100001100000011110100111101110111000100010011011111001100110000000100010001010101010100110000001111110001011111010000111100001111110000111111001101010001011111000000000000001111110000110100111111011100110100110001000011010101000011010011110011000000010001011100000000000100001101010001010100000111011100011101110011110111000101011101010000110111010011011101000101010001010001110101000000000100000001000101011100000000010001110011111111110000110111110000110000000101110011010001110001111100000100000001000111000000110101001101010011110100010001000000010101110100000011110000011101001101001101000100001101110101010101010011011101000001010011001100110100111101000011011111110000111101011100110000000011010000010011010011000111001100110001,2048'b00110011110000001111111111000001000000000001010111000001010111111101110100001101110000001100010000110100110100000111000011111100000001001100000011110011000011010011011100111101011111010101000100000100000100001111011111010000010011111101110000000001000001000100110000000100110100110011010100010100000111110111010101010000000011111100110101010000011100011101011111000001011100000100001111001111110111000000001100000000001100001101000000010111001100010000001100010001111101000011000001000100110000000100000011110101000011000000000101001111000001001101000101010100000001110001010111111111000111000101000100000111011101111100000000000100000111111111011111110001000101011100000100010011110001010011010111010100110011010011010100010000000000011101111100110011000100000111110111010011011111001100001101110100111101011111000101110101000000011100000000001111110011011100010100110100001111001100110001010100010000010101000111010100110101110011000000110011111111001101000000010001000001000101110001000001000100111100001100000000000001000111010111110000111101110100000011000000010101111111110100001100001100000000111111001101010000010000001111110111000101000101000000001101011101010011110000000000111100111101110101001111110001010001010001010111111100001100000101000100010011111101000100001111111111001111110011111100011111000000010000111100110100110000110001001101000000000100010000001101001101000000000000110011000111000000001111001100010100000100110001010000110100111111000100000011010000110100110001000111000101010111010011010111010100011100000100000001110000011101111111000101110101111101000100110100000111000100001101010000110101001100110001110001111111110011010000111100000011110100111100000000011111000100000000000011010000110001000100000101010100110100000011010100000100001101010011011111111101111100001101000000010001011100111101010111110000000000000011111111000011110000110000110001110101110000011111010011011100111111000111110001010100110000000100000000111111000000110101000011010001010111110101001101110000000101000001010111110100000000011100110000,2048'b11111101000000010000011111000101000100000111000011010111110101110101001111000011011111111101011111000000110000010101010000000000000101011100010111001111010111111100001100111111111111000000000101110001000100000100010011010001010100110011000000110000110000000000011100110111000100111111000011110001001111000011111100000100010000010111110011011100011111010101001101111101000111000111010111011100001111010000000001000000010011010011000101000000110011010111110011010011010011110001011100010101111100010001110111001111000001111111000000011100000011000111010000000101010101001100000100010000001111010011001100011100000111011111110001000111011100000000000000000000000100110011000101110101010011010011110000111100010100010101010001001100000011110000000101110001010011010101110000010100010100110000001100110001000001010111000101110111011100110011001100110000000011001111110100010000010111000011110001111100001111010001110001110011000111110100110000000001011101000101010111000000000001010101110000110000110000111101001101000101110111110000000000001100110100110001110000010011011100011111110000111100110111110011010011000100010011000000110000111111000101110011000011000111011100010100010001011100010000011111000000011111001101000000000011110101011111010111110101001101011111001111110001001100110011010011110001010000010001001100111111000000111101010000000000000111010000110000110101001111110111110011010101110011001100000001000111111100010011010101010011001101001100000000011111000000110000110001110000111111000111000000111101110100001100001101110101010111010100000000010101111111000111010100010011001100110100000011110100110000001100000100010101001100010000110111110011010011110101010001011100010011010100110101000001011111010111010001000101001101110001110011000011110111000111110011000001110000010111010000010011110011010011111100000101110001011100000100000000000001110000111111000001000000010000001111001101111111000101000100010011011100010101010111110000001111000011010000000000110101000101000111011101000001111101001100111111010100010000010001111100000001,2048'b01001111110100010100111101010000000111001100110011110001110000000000010000110011110101110000111101111101110111010100001100000000000000011101000011000111000001010101110100110100000101000011110011000100111111011111111101010000111111010100010100010011010100001101000000000101111111111100111111010101001100011101010101000100010000001101001100000001110011000001000111010100011100111100110001000011010000001100010100010011010111010111001101001101011101010011001111110001010011010101000001110100000101000101110100010100110011010100010000111100010100110111000100001100001111000000111100000000001100011101000100111100001111000011000100111101000100001100000000000111000011000000110000010000010000001111010011000001010100000000110001110001010001001111010100001111110000111101110001010001110001111111010000001111110100110011000100001100010011010000010011011101111100000000110011110001010100010000000000011100001100000000110001010000111111010011010100000001000001001101111101110011000111010100001111000000010001111100000100110000010011111111000111111111010000110111010100110001000011000001011111001100000111011100111101000101010001000100110011000011110000000100010000010101110100110100111111000000010100000100010111110011000101000001011101010101001100001100110100000111010001010111110111001111011100000011001111000111010100110001000100010001111111000100000000010101010101010101010100110000110101001111000001110111010101110001001101000111111101110100001100000000011111010011001101000011000000000000000001000000001101110111010111000011001100000001110011000111000001110101000011000001110111011101001111000101011101110000001101111111001100110011110101011101110101000000110001010000000001000111111111001100111100110001011101111111010100000111110000000101110101111111010000000011010001010111000100111100000001010100110000000000011100110001000000010111111111111100001111110101010001111111000000001100010000110001001101010111000101111100000100010011000000110011001111001101010100011101010000010100011101010100000101010011110001110100001101000011010011011111010111001101,2048'b00010100001111011100011111000100010111000100011100011100011100110001010100110000010011000001010000110001010011010000110001011100010001010011111100001100110111011100111100110100110100000101000111010111001111001101110011010000111101001100010100001100110100010001000011001100110101110011011101001101000000011100000001110101001101010011110011010001110101110101110101000000000001001100000111000001010111010011110111010001010001010101010100111101010101110101000000001100110101111111010011000001010111111101110000010000001111010011110100011101000001011100110101111111010001110111010001010001011100111100111101000100011111010100000001011111010001010111001111110100001100010011010101010001000101111111110000011111001100000011110011001100000000111100010001000101111100010100000000010000000011000001000011000000000101111101000100110011001111001111000000001100000001110011010011110100010100110111001111001100110001010100011111000101111111110100011100110000110101000101010111000000001101110001111100001100001101001111110011010100010111000001000001111100000101010011000011110011010000110000110001010011000001000101000000110000010000010000010100110100000111000001111100010111111111010100110001000000111101000101110011010011000101000100010100000100010101111111000000000000000101110001010100001100010101110101010111011100010001111101010001010001000011010101010100111111010111010011110000010000111100000000010001110100011100011101011111010011110000010000110101110001001101000101110000000000000001111101000000000011110000110100000000011111110111110011000000010111110000110000000101010001000100010011000101011100000001110011110101000000111100110000111100001100010000110101111100110111011100000001000000001111000111110101010001111101010111110100010011001100111100010001011101110011000111000001111100010011010001110000111100001111001100111111010000010001000001010101010011000001010011011100000111001111010101110000010100111111111111010100110100110100001101000011010100000001010111010000001101000000010011001101001100010001000100001100010001010000010001000100110001010100,2048'b11010100110000010101011100011100110100010000000100010100110001000000111100011101110100010101000100000000010100000101000111001111010100001100000111111100110000011100111101011100110101010101010000000101111101110111001111110101110111010011000011001100111111110111010100010111000111000101000101010111001101010000001100111101000101010000000011011111110111001101001100010111110000110001000111010111010111110001110001000001010001000101000100110100110101110100111100010111010111000000001111001111000011110111010111001111001100000111000111010011000001000111001100010000110100010001111111010100001100000011110111010000000011111100001111000100111100110011010111110011000000000111010001001111001101110011001101010011110000010000000100111100010001001100010001011100000011000111011100010100001101000101000001010111001101000100110000011111001100110100010001111101110111011111010001010011010000000001111101110101010011010101011111110011000001000111010111000100000001001111010111000101010100000000010011110111010000110000000011110000000001000100010000010000010000011111110001000000111100001101110011110000001111000000111111011100000011110000001100111100110100110111110111110011001100000001000101000101010100001111000000110000110000001100110101000111111111111101010000010011000000000101010000010000111111001100010101111101010100110100111100000001000011110011010111110111010100010000001100010100001111000111110001000100000000000111110111010111001111010011000000111111010100111100000001001101001101001100000100000001000000000011011111000100010111110000110111010000110001110011001111000101011100110000010101010100000011000100011100111101110011111101110011110011111111111111010101000000000100110111010111110000110001000000110001000011110011110100000011011100010011111100011111110100010000000001010011011111110111011101010011011111011111111101000100111100010100011111010000000001110101110100000001110000000101110000011101011101111100010001000100011100000111000101011100000001010101001100000101000000000111110000000000001100000101010111110001111111000111001111010111000001,2048'b00110000111101111101111111110001011111011111110011000001011111110100010101000111010100000100110100010101000100010100010011010111000000110100011101000000011100010011011111001100110100110011011100111111010111010000110000001100110111011100110100010101110100000100010101000000010001011100111111010011110100010001110000010000000111000011011100010001010011000000001101010000000111010011001101001100011111000000011101010001001100001100010011110001001111110000011111010000110111000011000000110111011100000111010100000011001111110011111111111101010101110001001101011100011101000111010001000100001111011100111100000000000100001111010100001101000001111100010100000111010000110011010011000101010001001101000000011100111100000100001111001101000011111100010111000000110011010001110011010011110001000111110111011100011111001111011100010011010101001111000000001111010100001101111100001111000100110000000011010101000001010000000011011111010001010001000000111111000000010001010001011111001100011101110000001100111111000100001111001101110000010011000101110101110100110011111100110100000000000111110111000111010001000001000001010111010000010101000101010011001111110111111101110100001100011111110000010011010001010000110111000111010000000111110001010101010011110100000101110100010001001101110100111100110001010101110000001100110100110001110000000011000100000111010100000011010001000100000000000000010111110101010111011100010100010011011101000000011101000001110000110000000000000001110111010101010000110011010000010101010100001101010001110001010101001101111100010011010100110011010101000000111101000001110011010000000101111100000000010111001101110001111111110001111111000100011111111101010111010101110101000000110101000011000011110001000100111100000100000001000001110011110111000000010011010100111100010111000001001111010100000001000111001111000001010001110101010100000100001101001101010101000001110111001100010100000001000001001101110100000001010101000001010000001111011101010100110111111100110100010001111111010100111111001100000011000011001100111101010111000011000001,2048'b11110001010100000100011100010011000101000101000000110000001111110111010000010111000111000011111101000101010001111111110111110011111111111100000100010011001100001111010011010001111100111100010101010000110111010001000101110001001100011101000101010100000001010111111100011101001101110111111101010000001111001111000000000101010100000111110000110000010111111100110111011100000101111101010100110000000100110011001100010000001101010001000100110011010000111100010100110001110101000000001101000011010000010101111100010011111100000101000011000000111101011101011100111111110111011101111100000011010111111111011111110101000100000100010100010000010000010101000111110111010111001100010000001100000101010001110011111101000011000000011111010111110100111101010011001100001101001101110001110101110011000101000011110001000001011111111111001111000111000100000101001100010000111101000001000001001111011100110111010000000100111111001100110011011101000100110000010001010111001111001111000000000111000011000101010001110000111111110100000000000000000011001100010111011101001100011100001111010000000001001111000100110000000000110111111111111100011100001111010011010101011100010100111101000001001101010111010101000011110001011100000100011100001100010011010001011111011100110000010000111111011101000111110111010001000111000100010001001100001101001111000001001101110000010001010100000001010100000100110000110100000111000101000101000011010001110000110101001101011101000111000000010100000100010111000001010001110001010111000001010011110011010011000101000000000011000000000000001101000001000100000000010011000001000100000101001111111100010001110100001101000100000000000000000101010000111100001100110100000001111101010011110000110111001100011111001101000001000111010000011101010000001101111111000001110011110001110001010111110011011100000001011101110100000111010101001100010100111100110111000001000011010100011101011100001111000100010000000000000011011100010000011100111100111100001111000101110101110101111100000101010001011100111100010000110100000001001101010011111100110001110011,2048'b01110000000000000111010000110101110000000001111101000101110011010000111111010100000101011111000100111101010000111111111111110011010011110000010011000001010111001100000111110111000101010000001100000100000001001111110111010011000000011101000011000000011100110101110011110100110000001100111101000100111111001111010001110100000111010001010100111111001101010001010100011111000000110001010001110000110011000101011100000100110100000011000111000001001111000000000100001101000111011100011101010111111111000011001100000100110001110101000111001111111111110011110101000111011101000111010111010001000100110100000011000100010011110101011100000111000001111111110111111101000001010001110000000011000100000011110101110111110011000001111101111100001100111111110011111101110000000000000011110001001100001111000000000000010111010111110000001100010100110001000101000001011111111100010011000000111111110001111101001100001100111111010101111101010000110101010100010011001101011111010111011101111111011111000000010111110011010000000001000000110101110011010011000100110011111111010111000000110001000011000000000011000000011101000001000001000111011101111100000001110011000100010101000000110111111100110011010011010100001101000111010100010111001111010000110000011111011111000100110011010111001111110100000000010101110000011100111111000011001111000100011101010101000000000100010100010100011100111100110100010100000011010000010011010100111101000101010000000011001100111101110101010101000100110001001101000011010011110000010000011111010000110011010000010100110011010000001100001101001111000101010011111111011100001111110111010100010111000011000111001111010001000011001100010011011111000001111101110101110100000100010000001111000100010001000101110100110100010011010011111111010000000001111111000000110100111100000011110101010111000011011101000100010011001100110001111101110111011111110100110000001101010101000100111101110011001101000000000100010011010001011111011111000100000001010111000111001100010001110100000100010101001101000101111111111111010111011100000100000111011111001111,2048'b01011101110000010000010100011100000111110001111111000101111100110100001111111100111111011100000001001111001101010011011111001100000000111111010011001100000100010100110100011101000101001111000011011101001101001100000001010011001100111101001101110111010001010011010111000011000001011100011101011111011101010000110111000100001100110000011100010000010001111111110101111100011101000100010000000111110011000000110000000000110011110011110100000111110001110100110101000011011100000111111100110011011111000101110001010100111100001101011100010001011111111100110001110101000100001111000000010011000000000001111100110111010100110101010001000011001100011111110101001101000111110100011101110111000111010011000000011101010000110001110100000011111111110011000000010100110000010000111100110101110001110111010100001111000011010001000111001100011100000111000101111100010100011101011111000011000100010100000001011111000100001100001111000101110111010101110011000111110111000001111111001101111111000100000101110000010111000000001101001111011101110111111101010001010101001100000100111111110011010111010011011100000001010111110011000000001100000100000000001101111100010111000001010000110000001100110011010101010000000011001100010000010001000100110100110101000011000100001111110011001111010101000111011100111101110001000101110111110000001100111100001100110101010000000011010011111100011111000000001111110000000000111100000111001100011100010000110001001111011111000011000100110000010000110000111100011100000000111100110100110001111100011101110100000011011111000001000011111101010000010111000000010001010011110101110000000000010111010000110001110101110001010011011111001111000101010000010001011100010101000001010111011100000100011100010000011100011100010000000111010100000100001111000000000011000101011100110111000011010001011111111111000101110001000111111100110011010000110111110111110111000111000011000100000011010011000100010011110011110001110111000101011101110000000101001101010100011100001101110000001100000001000100001111010000011101010011000001000001110101001101000000,2048'b00010011010011110100010101010100000000010101000100110011110001010011010100110000110101011101000011000101110111011101110001110100010011110101011101110011000100000111011101110001000101000000011101010011000001000000001101110000111111000011011100111111011101000011110011110000110101001100000000010000001101000000000001010001000100110101010111000011011100000011000111000011111111110011011111000011000011000000010101010000011111000001000011010001111101111100000011010100110000000101010000001100110011110000110001010100110000110100000000110101000001010101111111111100010111000100010011011101110001000100000101000100000011000000110100011111010111110100010101110000001100111101001101001100111100010000000000110101110000000000001101110011010000110000000001000011000101000100111111010111110000001100000100001111110100010011011111111101110000000100110001001100011111001100010111010100000001000101010101001111000111111100000100011101001101010001000011110001110000000100001100010011110011111111110000000100000000000011110000000000110000010011110001000101001100110101000101010000000000001101010011111100111111110101110001110011111111111111110100010011000100000000000101111111010000001111111111010111110111011100011101000111000000011111010000111111111100000011011101110101111111010000111101000111111100011100010101111111010101000111010101001111110000000101010111000001110001110011110100000011111100001100000101010000110100010001010011000001010100000111000001000001001100010100001100111101111101000100000111010100110011110011001100110000000011110111000011000111110001000011000100010000001100111111001111110001110111000111000011000011000111000100110111111100010000001100010001011111010001000011010011111100000111110011010011000100111100010101010000110011010111000000011111111101110100000011111101110001000000011101000000000101010111010101001100110001111101000111001101001111010100110111110101110001110100001111010100111101011100010101000101001101110011000101010101000011010001011100000000010000111111010100111101010000011101010011111100010100110001110011010011001111,2048'b00010101010101010101000001111100110111010001010000011111010000010000000001000011001100000000111111001111010101000000011101010111011100010011000100011111010000111101110101011111110100111101110101010000010011111101110011111111010011110100010101111111000101111100110000000000010011110000110100110101001101010000000001111111110000111100110001001101000111010011110000110000010100000001110000110111001100110011110001000100000101001101010000111100110001011111010100111101000000110000000000010001111101001101010111111111001101011100001111000000110101000000010011001100111101000011010000111101010011111100000101000100000101000101010000010111011101000001001111010100001101110000001111110001010111011100010000010001110101110101111101110011010000001101111111000000001100000100111111110111110001011111110000110000111100010111110001110101010101110101110011010111000100110000011100011101110011011101000011010100110000010011000001110101000100111100000111001100011100000011011100011100000000010111000000110000001101110101110011110000110100011111000001011101000100010001110000010101000011001101010111000100000011110000111101000100010100111101010101110011001111110100010101010101110001110011010011000011111101010000000111011100110000110100000111010100000001010100110000010001110101000011111100111111010001000111111111010101010001110100001101001100010111111101010001011111011101001100000001110011000000110000111111111101010100000111000111110100110011011111011111111101000000110101110001110100001101000101111100110011001100000111001100010101011100001100010011001111011100110100000011001111011101110100010000000011110100110001110101011111000001001100010100001100111100110001010111001100000100000100010101001100110001010000110101000101110100110000110011000011010101110000011101000111000101111100110101010000010011000011110001010000010001111101110011110001111111010001110111011100001101011100010001110000010011001111000000000000000101010000000100011100010011110111011101000100111100111111110011110100010100010011010100011111000101111101000011110101000001110100110101010100,2048'b00010001010001000000000011011101010011011111110001001111011100000000111111010011010101000011000001010101110100000000110011000001110100001100110000111100000000110000010001001100111111010100000101111100010100010011111100110101000000000000111111011100000011110111001101110100010000000000001100000000111101111100010101010000010100110101000001110011010101010111010000111100000000000001001101010101000011010011000000111111111101010011110101000011110011000000010101110000000001000001010000110100111101010001001111010100001100010101111111000111111100011100110001000111010100000011010101000101000111111111000011110000010100110101110000110100011100110001010111000001111100000100110000010100000100110000111101110001001111000011000001001100111111011100001111011100111101111100001101001101110001010011000111000111010011001100000100111100110000010101000100011101000011000000010101000000010101010001001111010100010111000011001100111100010101000011010000000000000001010011110000010100111100000101110000000101011100000101000001001111011100110100110111010111000011110001010000010100001100000011110001011100000000011111000100110100110101010111000101000000010100110000010001010000111100110001000101000011000100110100001100010100000111000011010111011100110000010011110000110100011101000000111101111100110101000001000001011111111100110100111101111100010111010111010101000000011111010100110000010011110000000111010111011101011101110100001101010100110101001111110011110011111100011101111111111111001111011100000011000011000101000100111111111100011101110101110100011100001100000001010000110100110101000111110101110111000100001101001101000001010001010111110000010001010100010001111100111100110001110101000100111111000001010011110011010001111100110000011111010111000000011111011111010100000101001101000001010111110001001101000001010100110001000100001100001100011111000111000001110001000000111100001100110111110100110001111100010111110001010101001100000111111100011111000001110011110101010100111111110100111100110001000011000101001101000000010101000000110101110000010101110001,2048'b11000000110101111111110011110011000100000100111101011100000000000100010111011100010001110101001100010001011100110101011111001100000000111101001111010111001111000111001111110100010011011100010011010111001100001100000100001111010111011100010000001100000000010000110101000000111100000011110000000001000001010100010011010100110011111111001101110001010001010111110001000001000000001111001100110101111101000001001100000001001101001101010111010111110111001111011101000101000101111100110001010011010101000000000111001111000011010011001100110100010000000011110001001101010100000000000000000100111100010000111111110100000101000011000100110011110001000011000111011100010111001101011100010000001100010100010100011111011100011101010100000101000000111100000111110011110000001111000100001111110000110011010000001111000101001100010100011101000011010111000011011100000100000101011100110100111101000011000011000100001111010000010001110001010101110011110101001100110000000100000101110001111100001111000011001111110111000001110001110100110000010101110001010111001111011101000011010011110100110001110100001101110000110001000001010101110001110100011101010001110000111101110011010101000100110100000011000001010001010100011100000101000001000100000000000101011101110011000111110100000000110111110001110100000000001100000001111111111111010011110101110001011111011111010011110000001101000100110011001111110101111100000011011101010001010000011111010101011101000101010000000000111111010001001100001101010000001101000011110000111100111111010011010111111100010011010001010101011101000000010000111111001101000011000100111111011101001111110101001100000000111100110000001100001101001101001101011100110111110101111100010111001111010001001111000100000101011111000000110000011101000000010000010111011100010101000100110000111101010001001101010100001101010100010000110000110000110001000011000100010111001101000101010101111111010000010001010001110101011101000100110011111101110100001101111101000100000101000100000111011100110111110000010011010000000011010111110111010001010001010000010011,2048'b00001100000001010111010100000000000111010011010101110000011100000101000001010011000100000001001101000001110001110001001101110111011111110000110100010111110011010011110100011101010100011100110001110100010000000101011100110101011101011100010000110100000000000111000000110100110100010011010011000000110000000011011111111100001100011100010100010011010011000100010000111101001111011111011101110000000000010111000000110000011101000000000000000000000011110000001101001100010100010001111101110011000100111111010100010101001101110101010011010001010100000001001111010100110000111101001101011111110000000011000000010011110100011111000001010011000100111111010001111111001100001101000101010000010101010011010000110111000100110000111100111100110001110011000011000000010111000001110001011100110100001100001111000011110000001111000100010101010111010000000011111100110100001101000111010101110001001100001101000001110101110001110011011111011101000011110000010000110011001101000000111100011101111101000001001111010001111111001100010100110000001101000011011111010000000011110111000101010001001111110000010011000100111111000111001100000100110111110011000100110111000111111111010001110001010000000111000001011101010100110001000011010111010101000011110000010011001100111111000011010001001100001111000001010100010100000101110100011101000000010111110011110100001100001100000111000000110100000000010111110000110001000100010000110101000100010000010011110111000011001100010101110100110011001111001111000100000100010001011101110001000001110100011100000001000011000000001111000101000101001111010100010011000111000111000011110101010001010101110000110100001101110000011101001101000011010001110011110111000000000100001100001100011111001101111100110101110100000000111111001100110101011101000001010101001100011100010000001101111100000011000111110000011111011111110011110101110001111111111101111101110011001111010001000111011111010011011100111101010000111111000101010100001101000111000000000000110000001100011100000000000011111100110000001111001100111100000101110000110100110101110001,2048'b00000000010100000000010100000101111101111100110101011101000000110011110111111101000100000001110101000000010000011101001111111100001111001101111101110100111111010000110111111101000101000100010000000100000011001100111100010001010101000001110111010000010011010000000001110101000101011100110000001101011100000101010011001101110000001101010000010000010101010011000101010001110011110111000111000011011100010000110011010111010001000001110000110100111111110001001111000000111111110101010001010100000000111101011111110100110001001100001101000000011100000011000101000111110100011100000101000001000100000101010100001101110001001101110101000011110101110011111100001101010000111101110011010011010100011111010011000100111101010100111111010001110111010100111100001100010100011100000100011100001100110001010001110101001100110111010000000011001111000100000111001111010000000000010000010111110000111111110001011100110111010111001101111100010100000000010100000111110000001101111100010000011111000000111111001111010001010000110011111101111100010100000001110001010100111100010000111111000000010011001101001101000100000101010000010101010001001111010100110001001100010001001100000111010001110100010101000100000001010100000011110100001100010001001101000111010111001100000101010011010100111101000000110011000011010100111100010000000001000100000100000100000101001100010100011100010000000111000000000001110001110000111111011101010000000000110011011100000001110000000001000100000111000111011100010000110000000111111101011101011100000111001100010000110001110011110000010100010100110111110000001111110000111101110011010101010001001100001111000000111100111111000001110111001111110111001101011111110100001100000111110100110000010101001101110000111101010001110001001101010001010101110101110111110000001100010000000000000000110101110101110011000001010100110011011100010101111100010111011100000111010011111100000011110111010100000100110101011100000001001101111100000000000111110100011111010100000101011101111100111101000101000101001101001100001101000000110000110000110111110000000101,2048'b00111101000101000011010000000100010100000011110000110001000011110000010100110011110100000000011101000100000111001111000011001100000101110000110100001101000101001111010000001111000001110011011111110001001100011100001100000011000111110100111101110001110000111100010011000101010111001111010101011101111101001100000100011101010011001101001111000001000100000100111101010001110101001111110011000001001111001101010111000011000011000000111100110111000100110111111101010011011101000011010100001101110100000011010011110001000000110011110001001111010100110101110101110111000001110001110100001101000100001100001111000001000111000101110101110001010001000100000001111111001101111101010001000101110000000011000100011101001100110100110001011100000000110101000001010011000101000101111100000100010000110100010011110100010000010111010011000011010100001100011111000001110000000000001101110100010011110111110000111111011101110000111111110011010001000000111101110001110100001111010100001111010011010001001101110100000100000111110001001101110100110011010100010001000000000111110000011101110100000001000001010100110101011100001100000011111101000111111111111101010000111101010101010000011111010011010100001101010000010000010001011100111111111100010001010100010011110000110001110000110100110100000000011111110111111111000100010001000000010011001100111101010101000100000001110101110000110000011100000001110001110100001100010111110000110100000011000000010111001100110000001101000001110001001111000000011100000111001101001111010011110001001100111101000111000001110001011100110000010011110101010001001111010011001100110000111101001100011111000001111111000111110011110111000100111111001111010011010011110000111100110111010011111101010101110011000001001100001101110000000001000111001100111100001100000000000000000100001101110000010011001111111111010100110101000000000100010011000001011111010011111111110101111100000000010100001100010001110000010000000000110111110000010111000100011100011100010001110100001111111111110101001111110000001111110101000111011111000000110001011101000100,2048'b11010000110111000000110011010111110111000000110000110111010011011111011101001101010011000001110111001101001100110001110001000000110111110001000100111101110011011100010000110100110000010011110001110111010100110000110011011100001111010011001111110011011101000101110101000000000001010100110001010011000000110001010001000001000001000100110000000100000101000101110111111101000100110111000100111101001101010101110000000011111101001100110100011111010011001100110011110001010011000011000000000001110001010000011100010111110101000111010100010000010001000100010000110100001100111100000100110001011111010100000000001101000101010001010100110001000000011111010100000101000001000101001111110101110100001101000101000011000101001100000011001100000101010011010111110001110101010111001100110001010000001111010101001101110011000000110111110111110101010001110000110000011101110000000000001111001111011100110100111100000111111111011101011101000101011111000101011101000000000000110100011100010111000101010111110000000100111100110000010100010001000100010011010100000111000100000011110100110101000111000001011100011101111100110100010100010011010100000100110111000001010100010111011111010100110000000000001100000000000011010000010100111111011101001111010100110101110001010111001111000001010001010101011100110100000000110001110001110111000001000000010000010000001101110001111100001111000111000000111101001111110011000000110011010101110000110100011100111100010000110011000000000000010000000111111101010011110101000000000001010111010001110001010000111101010001001100010011011100111101011101000100010101001100110011010111010011001111000000110000000001010011001111000100001100010101000100111111000101010001010000000011000100001100111101011100010100000001010000001111001100110101111101000011110001010001111111111101001100110001001111111100010100000100010000010001011111011100000001010001010011000000001100000100111101000000111101011111011100110001010011000101011101001111010111110011000011011111010000011100010000000101000100000111111101000011110101110100010000111111010001011111,2048'b01111100001100010100110011010000011100000001111100010101110101110001010000000100110011011101000000110100110100011100110111010001010001110011000100001100010011001100000101001100111100010011010100110101110001001100111101010111001100110100000111010000000100110101010111000101010001010100000000110100111100111100111100001100000100110001011111010111001101010000010011010100011101010011110111010111110001110100110000010011000011011101110000000000110001110000011100000011001100110100010001010000000001011111000000011100000001110000000000001101111100011100110100011111110111010111110001010101000000111100111101110101010011011101000001000000111111010011000000010000111100000111110011111100000001000101011101000011000011010000010100001100010011111100000011000101010100000111010000110011010001000100110011000000111101000111000101110101010111000011011111010001000101011100001111010000010011000000111111000101011111110001110000000101110011001100111111000000000111010001111101001101011111011101010101000111111101001111111111010111011100001111110111000111111111110100110000110000000100110011000111110111010100000011110011001100010111000001001111110100000001000111010001010000010000110011001111011111010101010001000111000101010100111111011111010100001101110100110000110001010011110001011100111100110100001100000111110100000101110101000101010011011111000111111101000101001100011100001101110101000000011101010001111101111100010001000011110001000001000101000000010100111111001100000111000100010000010100110011110111011101000011010011110101000011110001110011110011000011001100000101000101000000110100010000110111110001110100000000000000000001110111111101000011000100111100000001000111000100001100010000110101001101111100010001011111011111111101000000000001010101010001000101110000000101110111001101110000111100010000111111110001011111110000111100110000111100000100111100001100111100110000000111111101000000110000110111001101010001110111111101011100001111110100010000001100111100010111010000001111110100110000011111011100110001011101000001001101011111011100001100000000,2048'b01001100000000010101110100011100110011010111111111010000000111000111010011010000001101001100110011011101111111001101110000000001110001110011111100000111001101110000111100001100010011000001000000110101000000011111010101000100110001000111000001110111000000000111010100011100011101000001110000111111110011000111000011110101010100011101110111010011111100001101000011110011110101000011000000110101011111000100110000001100001101110000000011000000011111110000110011000100000100000001001111110000011111000111110100000011010000001101110000000101000000010011111111001100110011011101010101111101111101000100001100111111001100110100010101001100111100011101000100001101000111011100000011110101010101011111010000111111010100011101011100110001010011011100001111110100010000000000000100000111110001111111010100111101001101010111011100010111110111000000010100011111011111111100000111000101111111000001000100110100111100010101011100110011010101000100011100001100010111110011010101010101110000110000000011001100010000110101111101110111110001000000110001110001011101111100010100010000011100010111001111000100111101011100011101001100011100010011000001111111010011000100110100111101010111001101000000010100110001110001000001000000000011111111001101110101001111001100110001010000001111110100110111110001000000011111110111000000000011001100000000010001010101110000000111010001110011111101010101001101111101110111110101000111111100000011110000011100110101000100000001110011110100011101010001000101110011000111110011011100001100011100111111000100011100010011110101000111010000110011000000010011000101001100010111000111011100010100110111000000010111001101000100111101000100010000110001110011110011011101001101110000010000011100001100111100010011010000110100010001010100010101010100110001000000111111110011110001011101000011110100110000000100000111000000001100000100111101110100010100011101010000001101000100010101110001110111110000011111110111010100000111000100110111110101000000000001000101010000000000000000000000010000110100000000000000011100000101001100000001010111010001,2048'b00111101011100000001110000111111011111111111000000110101000011110000010111001100110111000101110000001101110101001101110100010111000101010111011100110001110000010100110011010000111100000000110001000011011111110000011100110011000100111101000000011101110000011100010000010100111111000001001100000001110000011100111100001100010001011101001100011111000001011111000101000011000111111111000000110100000111010111110111001101010000001101001100010111111101011111001111010000001111110100000011110001110001000111011111110111010100000011111101110011110001110101000001111101010011011100000101010000001100000011000101000101010011010001110111000100110100001101010100000100000011011101000000001100010111110011000000111111010000010111000101110111110011011100110000010000000100010011110100000100001101000101000101000101000011111100010001000000001111000001110000000111000111001101000100110111001111110011000100010101001111111101000101110000010000000011001101011100000011011100110000001100010001111101000101000000010011010111111100111100011111110100010001000001110000010001111111001100011101001111000011110111001100000000000111110000010100110000111101111111000111000100011100010100000100010001010000000111110000000001110000010001000011001101011111010101110011110000110101010101010011001111111100011100010000001111001100011111011111110111000011010100011100111111111101000011000011000001010000110101010011010111011100000000110000000000110100010011011100000100110001110000111101010011110100011111110001000001010101011100110011001100010000110011001100011100000011011111000001000101010000111111001111111101000111110000011101011111001100111111000011010111000101000011110101110101110000000000110000110101111100110011001111010101011101110100010001000111110000001111110100001101010001110000110000000000111101110011011100010000010000010100000011110000010100010111010100111101001111000101011100000111000001001100010100000000000100001111000000000001000000010001010101000111110001000011111111010011111100010001111111010100010111001101000011111111010001000111001100001111000111111100,2048'b00010111110100110100110111001100000000000001001101110101000100000101110100011101110011001100011100010001111101111100010011110100010111001101000100000100110001001101010000000011000001010000001101110011001101010000010111011101010001000001110100000000011100000101011100110100000001110000110011011100001111000000000001000111000011010000000101110111110001110101010100001101000100010101000101110101111101000111001101110101001101010001000101000011010001011101000000000001110001010100110011000100010001110011010000000111011101000011010111111111010111110001010100010011000001000011001100000111001111110011001100010011000001000100011101110100011111110000000100110011000101010001001101011101110011011100010011000001110000000000111101110001110100011111000111001111010011111111111111000001000001110111010001011101110111111100010000000011010101010100000001000100010001001111001100110101010101011101011100000011010101110011011111000000000000110000010100010100000101000111010111010001110111000100000111111101010000110001000101000000110000010011110101010001000000010101110100000111011111110000010100001101000001111100011111001111010011001101000101110011000100011100010101011111000111010100110001011100111100011101011111001101001100000011000011000011110000111111011100000101010000000000110000000100110100001100000001000101111100010100000001000011011111000001010100010001001100000100001100010001010111001100010000000000000001110001010101000011011100000100110111000000011100000101001101011100010000000111111101001111000001001111000011010001111101110111010011110000000000000001010000111100001111010001010101001100111100111100111111010100110011110011000100110011010011110011010001011101010111010011011100000111011100011100011111110011000111000011001100010100110011000000110100010000011100011100110011000111110101001101111101010001000000010101000100111111010101110100011101010111011100000011010100000000001100110101001111110001010001000011010111110000000011110000000011111111000111001111110001110001000001010100000100111101110100111101010111110111110000010100011111110101,2048'b01000000110001000000010100110101110001001100011100010000001100110001001100110100001101000000010101111100111100000000010111011101110000110001111100010100110000010101110101000101000000001101110001110011000001111111011100110000010011000001010011001100001111000001001100010001110101111111001111010111111100110011011101011111010101001100001101110100000000110100000111000111010011011100000111010001110000010011000001011111000011010000111101110000110111000001000011110001000111110000110011000100111100010101001100111100001101010111110000010000000101011111110101000100010101010101000001011100111111000000110000001111001111001100000011111111000101000000000011110000001100010111001111000000000111110011000000000000011111010101110101110101000011000011000001110111110000000101000001001100111101110000110001000101001101110111000101010111001101001111001101111101000011001100010000011111000101001100111100110001000000001111000111000000010101011100110000000101111111110101110000111101000100010011111111001111110100011100001100011101010000011101001111010111010111010011000100111111011111010011111111111100010111000001000001010100000111000111010001000111000101111111000101001101111101110000000100010001000001011100000111110100010100011101001111000100010011110100110001001100110000110111001100001100111111110111111101110011000011110000010111000111001100011111001100110011011100001111000100110100110111110001010001010101010001000011110000111100010000011100000000001101001100010100001111000011010111110000010001000111110000110000110100000001010001010001111101111100010100011100000101001111110000010000010100111101010000010001011111010100000011010111001100011101111100110011111111000100010000010100010100010111110001011101111101110001000011110011001100110000000000011111000111110011110000110011000111110000011100001100000000001111000011011101111111110000000011010000110000000001001111110011000001010101000011010000110101000001001111000100110111000001110111000100010111001111001111010011000001111100110011110000000011000011011111111111011101000011011100010011000011110011,2048'b00011101111101010011001111011101011100000111010011000011011101010000010000010101010101010101011101001100001111110101000001110000011101111100011100010000000111110100000101010000111101000101000011111101000000010101111101000011110000010100000001110011011101000111001100110000000100011100010101000011110111110111010011010001011100110000011111010101011101001101000100000001110101010000000100000111010000110011011111000100110111010001000111000101010000011100110111111100011100110001110011001100010100000001000000010001010000111111000011000100000000000011111111110100010111001111000111110000000011000111000100010011111100110100010000000011110000111100010000000000011100010001000100000011001111110011000000111100110011010011111101011101110001010100011111111100000000000100000000110001001100111101010001000111010101000101000000111100110000010100111101000011110100010001011101011111010001010001011111010000011100000101111111001101010111001111000001010000000100110000010000011101110100000100000000000000000011111100110100110111000000010001010111000000110101010000010100000000110001000011110100000001011100110011011111111100010011011101001101000100111100111100011101010100001100000101011101110101000101000001001111111100010001110000110100011111010000001111110101111100010111010011000011000111001100011100010101000000011101000100010001000100010100110000010011000000000100110001000100110100001111010111110111010111001101010100000100011101110000011101000100010111000001110011001100010011001101010001000101111101001101010101011100110101010111000101011100011111010001000011001111001111110100000011011111111101110111001100110101111100001101110000110101110001010001010100110000000100010000111100000100000001010011110100111101000000110100110001110011000011000011001100111101111111011111110001010011111101000000000111010001011111000111110011001111000011010011010011110101011101000111010101000100110001010111110001110111000100111111001111010001000011010011110100000000110101000100010000000111110001010000110011011100000101010011010001010001000101111100110000011101010001,2048'b01010001110000011100000011001100010001010001110101010000000101011100010001001100010001010011000001010000110100000111110001010011110111000000010011110111000000011101011111000100111101110001000100110111000011110101000000011100000011010111110000110000010101010111000101110011000100110101110100000011110100000111111111111100110001000111110000001100110101000001110101010000111111110111000101110001110101001100000111001100010100010100111100110000110111000100001100000011010011010101010111011100111111111111000100010011011101001100001100111101000001000000001100001101110001011100010000001100110001000011011101110011110111001100010111111101000111010001011101011100000100000100111101001101010011010100111100011111011100000011110000000001001100110011001100000000110111000111000000111100000001011100000000000001001111010000111111110001111101110100010000110001010100000101110100011100110100000000110001110001110100110101111100010011110011010000110111110100000101000100000100000011110000000001000101000000010111001100111111000000000000000011011100001100010001010011010011000011000000001111110100010000010001001100000001010101000101110100110001001100001100010011110000010001000111010111110101001100010001010011110100111101001111110001110111000100000001111111011101001100110011010011000111010101110001000000010100001111110000001100110111001101001101010000001101000101010001010011001111011100001100110011010100010011110101010000010101000000000011000100010101000111111111110000110011000100110000000111000000000011000011001100010101110000110100001100000101010001011111110001000000000100000101010101011101111101011101111101000111010011000100010101011100011100111100010100110000000011000001110100000011010101000100000101110111000000000000010100010000001100010101000001001111111100010101010101010100000101001100110011111101111100111111110000110111001111010000001101110011000101110011110011000111110101000000111100110001001101000011000011010011110000011111110000000001111101010101110000010100010001000000001111110001110011000000010101011100000001010000001100000011010100,2048'b00000000110001000011000101000001000000110011111111011111000100001101110000000111000001000101010100001101000101110001010000001101111100000101001100011100010001000101010001111100000001000001111101000011011111001101000000010000111100001111110111000001000001001101000001010011110100000101001100001111011101000001110100000101010001010111011100110101010011001100011101010111001100010100110011110011010001010101010000001111011111010101010101000000111111001111110001110111010000011101000101000000010000001100010001010100010101110100110000010101111111110011010100111100000000110000001100011100000000010000011100110101000101000100110000110001110011001100010100010100011111110000000011010011000011010001110111000111010011010111010101000101010100110000000100010111000000110011010001000000000000011101010011001101010011011101010111110101010101011100110000001111000100010001000111110101010100000001001100110000110100011101011100010100001100111101010101111111110111110100111111001101110101000101011101110001111111001101011111000001010101110001010000011111111100001101000000010001000111000100000000001100110000110000010100011111001101001111011100011101010000111101111100010101010000000001111111010100000111000101110100001100011101001101011101110000010000011111000111111101111100011111110000000011111101001100110011010100110101110100111111110011001101111100010011010111000001011100110111001100010000000001110101000000110011010111111100001111000100010100110100000001110100110011000111011100010000110000110000010101010101000000110100000000110101110100111101110100000011110000110011010001110100001111001101110100110001010001000011111111000111000001000000010001110011000001110101000001110111110111010101000101001101011100000111111100000100110001011111000011000011111101111101000011110100001111000011000000110001110001001101010111001100000011010100111111010101001100000100000101001101110001000100111100111111000011110001111111001111000000010101010011010100111101110011000001001101011100000100001100010011000001010100011100110100000100010000110001001101010101000000111111,2048'b00000011001101010101010100001100010001000101000101000001110011000011110001110000000000001111001111010101000000010011011101000111010001110001110111011111110100010111111101000101111100000111111101001101010001111101110001110011111100110100000111111111110100010101111101010000000100010000011100000001110011011111000011110000011101001111011101010111110001000011000111010001001111000101000000110111110100110000001101000100000100110011000001010100000101111101110000001100110001110000111100000001000011011111010000110111011101001101111100111111000111110111110001001100010100000011000001110011110101111100111100000000010111000111000000010111110011011111001101000111000100110011000101000011011101000000010101001111000111000001111101010011000100111111010000110100010100110001000111010001111111001100110111110001000101010000010100010011010111000111000001110000010111110001110011110111001100000000000000001100000100110011011100000100110011010111001101010011001101010100110011111101010100010000000111001100000011010000110000001100000000000011110111010111001111110100111111010101010001000101010011010101001111001100111111110100110111110100010001010000001101010100000111111101001100110001010101110011010011001111010000000000000011011100110000010000110000110001111101110101110100110101110001110111010000010111000011111100000001000001110100000000011100000000011100010001000101000101000000011111000101110111000100000000110000010011010011110100110101000001000001010101001111010101000001010100001101010000000001010100000111110000000000010000010000110000110000111101011101010001011101001100000011001100111111011111110000110001000100010100000001001111010100000011011111110011000011010111010101110100111111011101111111001101110000111111110000000101110001000100001101111111110011000000010001000100010000110001111101010011000111000011111111111101000101001100110111110000000001000101010000000111010101110111000100000011011101010101010111001111010100001111011101010000000001001101111100000000000111010000000100000001000111011101001111110100001111110001000011011100110101110111,2048'b11111111011101110100000100000100000011110011110011011101000000111100010111000000001111001100010100111111000111010100011101110000001101110000011101111111001100111111010101001100000100000000011111110100111101110011110001011111110011001101110101110101111100001101000000111100110000000000110101010101000101000111110100000000000111110101011101110111000000110011010000110111000011001101000000110101110000000000010101010100010101110000110111110101001111000111110000110001111100010001010101010111000000110001000000110001000001000100110000000001001101000001000001110001000001000001001100110011010101011101111111001101001100001101111100110001110001000000110001001100000001110101110111010000010101010001010011110111000001110000110111110101010011010100010001000100010000000011111111000000000100000111000101000000111100011100110001001101011101010001000101010000010100011100000011110000000111011111111100110011010001110100000011010011110000000101000101110001110111110001001100111100000100000111000101000101001101110001001101000100000111001101110111010101010101000011011111111100110111000111001111110011110001010011000011111111000000000000010111000011011101110001110101111100111111000101010000010011110100000000000101000000000001000111010101110101000000111100010001110111000111110000010101000101111101011101010101000111010111001100110000110001010001000100010100111111010011010011111111111101001111001100110111111111011111110100011100010001110000001100001100110101001101001111001101111111001100000101000101010001000000001100001100000000110111010001110101001101111101010111111111001100111101110000111100000101010001111100010101011100000000000111010011110111000000010011110101000101000000000001010001000111010111110011001111000111010000000001000100110011011100001100010001111100000111000101000001010000110101110011001111110101010100000100010001011101010000000000000001001100010100000000111101010111110000010001011100000100010000111101000101001101001111001111000001000101001111010000010001011100110111000100110000000000010111000100110111010001001100011101000101010011,2048'b11000101001111011111000100110011011101000111010100110000010000110000110011000001010101011100000000110101110000011101000111010111000100001100110011000100001101111100011100010100001111000111000111011101110000110011001111000000010100010101110001111101011101000011010000010011010000011100000001111101110001000111010001110000111101111100010000001100000100110000000001000011000101110000010100010100110011000001000100011111010100000101111100000100110100010100111100010111000000011101000100000000010011000001000100011100000001110000111111110011110100110100000101011111111100010011000001000111011100001111000011010100000001010001110000110000010001110001110011111100110011010011000111110100000000110100010111000000010111111100000100011101110000110000000000010100010000000011011100000000000011011111000001110000111100010001010101110100011100010100110111001111000000010100111100010101111101110001000011000111000001001101011111000011001111110111010111011101000111110001000001010101000000000000010100010101110000001111010011111101000001000100001111000011000000010100010001000001010100001111010111010100110101010001001100011101010011110011111111110001110111000111000000000100000000000100110011010100110011010101110101110111000001110001001111000011000000000101010100010100011101010111000000110011000000000111000011000001010000010011111100000001110100010101011101010011011100110001011111010000001111000001011100011100010100000111001100011101001100111101111111000001110100111100011100010001111101000011110100000101110011111101110000110111111101010100111100000001010000011101010000010101110001001111000111110111001101010000111101000100010000010000011101110001110000110001110111111100110101010001111111010001010001010011110011001100010000000100000100010000010000011101010111000011000000010001000011010100110000010000010001000101110101010001110001000101000000000001000100000000110101110011000000010011111101010001110001000101000011000100000001001111000100000011001100110000111100000111110111011111001111000000000000110011110011110000000100000101010101011100010111011111,2048'b01010011110000110100000111110001110000010000000100011100001111010101000100110011011100111100010100010111000001110011000101110000001111011101111100000111110000001100000100001100000001010101011101110111000000010100110100011111010000000011000000000111110111011111010001000001010001000111000111110011000011010011110101010111111100010000000111010001010000111100011111110111010111111101110100000001000100110001000111110001001101111100110000001101011100011101000101110111011111000100111100111101001101010001010000010011000011000000001100110000010101110001010100010011110000010001011100011101000001000000011100110011001111010100110111000111000000111101000011001101000011111101000101110000000011111111110100010101001100000011110101000101011101011100000101110001110101000000111101010000011101111111010100011111110100111101110001110101110000011100110111001101001101000111110000010000111111011101001111000000000011110100110001110011111100001111001100000011010101111100110011111101010011111101000101011100000000000011000001010011110011111111110101011100010111010000011101001101111100010011110001000100110001001111011100010111001101000111000100000000010100110011001101001100110100011111010011001100000111111100111101001100110001110000001100110111010000110001111101001101110001001100110100010011000101011100110011110111001101110001011100110011000101000001010000001101000100011101010000001100000011110000000000110100111111110011110000010111001111000000000111011111010100010101000111110101110011010011010001110111111101010000110111001111011100001101110000000000110011111101010111010100001101110101110000010100111111010000010101000100111101010011010100011100000011011100000000110111001100111100110011110011000001000111000100000111010011110001110001111100011100010011111101000000010111000001111100111111011101111101000000010000110100010111011111010111010111110101010011010001110000010000111101111100000100010000000001010100110111000100011101011101111111000101011100111101010111000000110000110100001100000001001101000000000101001100000101010100110011011101000001110011,2048'b00110101000001111101000001011101110000000100111101001100010100110001000000111100011100000011010111000111111111111100010000010000110111010000110101111101000000000101000011010001001111010000001100010000000101110001010001010000010101000101000000110111001101010001110001010011010000011101111101110001010100000000110001110101010011110000000101000111000000001111110001000001001100111101000100011101011100110000011100001101110000001100111100011100000011001100000101110111001101010111001111000000011111110111010000011111000101011100110100000001010111111111001111010001111111001101000000011101001111000011000001010101000100010101010111000111000011001101110001111101110100010100111100110011000000010100000000010000110000000001000001000100011100000001000100110011110101000000011101011111011101010100010101010001110111000011010001000100110001110011110001000011010111011101111100001101000001011101110100010100000000110011110001000001111100110000000011110100001100000001010101110100110000110000011111010000010100001101111101111111010100000101011111001100000000000100001100010011010100000100110100011100110100010100000111110100001100000101111111000001110111110011011111000100010101000100010101010100001101000101010101010111110011010100000100000001111101000101011101110001000000000000111100001100000001110000001101110101011111111101111100000111110100110111010111000001010000010001011101110001011111000100000111110111110011010001011100000100000000110111110100000111111100111111110100010101110000010111001100110100110011111100010011000111000000000001000000110011001101010101001101001100110000010000110001000111110000010000000100001100110001011100000101110000110100110100111111110101111111011111110000110011111111011100110100110111000000110000110011000100011111111100011100110000111100110111000011110011001111010111110011111101001101011100000101110011000011001111111111010101000000001100001111110000111100011100000001010000000001011101010101011101110001000011110100111100001100001101000000110101010011110100000100001111000101010011110000000011110101110100011100111111,2048'b11111111001101110011010111110111001101000000000001010011000000011100001101010001000101001101000000000100010111110000000000110100111101010101001100001100000011000011010011001111111101011100011101010011000100000000010000000000001100010100011100110101110100010011010001110111001111011100010100111100111101010001010011010001111111011100010100001100110111110000111111010011010000110100111111111101010011110001110100010011000100000011111111110000011111110000000111111100000011111100111101111111011101000100000111110101000100010101001100010100001100110111000100000111010000011111001100000101001111001100000000011101110111111111011111010100001111010000001101011111011100010111011100010000110101110111010011000001110111000001010001111111110100000001011100000100000101001100000101010101011100010100010001010111010000000001000011010000110000110001110111110000111111000001001111010100010011000100001111110011010011000011010001010111010111110000010001010111011101110001111100110011000001000011010100011101010100110100001101110100010011001111010111110000010011000000000100000000110111000111110001110000110001111100000101011101010011001100010000010011111111000111000011110001000001000101000000110111010101000100011100000000001111000111010001000000110001001101001100010011010100010011001101000100000011001100011111010001111101011100000011110001110001011100000111010000011101011100110000010100110111010001111100000100010001110001010000011100111101010001011100000011110111110111001101001100000000010100110100011111001111000100110000010101111111000000111111111101000001011111010000110100110101001111000011010111110101111100000001110001010001111111110111010101000111010011000111001100001100111101011111000111010111001100010011010001011101000011000100000011110111000001001100110001000011010101111101000111000011110011001100011111000111001100001111000100001100001101111101010011010001110111001111010001111111000000000101000000011101111100001101010000001101010011000101010100010101001111110100000100000000011101000101011101000111010000000111110011010111001100001111000000,2048'b00110000110111000011000111011100110100110101001100110011000000110101010101110111110101000111110011000101000000111100110100010000000000000100000011110001110111010101000100010001010011000100111100010000000011000111110100011111000001010011110100010000010101011111000001110011001100110101010100010011111100001100011100010000001100111111010101000011010100011100110100000000000111110000001111110011110111001100010011111111110001110111010101000101000011011100110101010111111100011100000001010000000000111100000100001101000000110000010001000100110111000001001100011111000011000011011100000001110100000001110011110000000000000100010011000001110111010011000101000101011100111111000011011101010000110000010101111101110111000001000001000000001101001101110011111111010000001101000000001101010111010100001100110001000001110000110100110001000001011101110100010000010011111111110111000011110011001101011100011100111100110100000111111100000000110100011101010001110011010101010101010111001100110001110011111111001101000111110100001100001101000111000000010001110100000001000001010000010011111101110000011111110001010001001101010011000100000101011100010011010101001111110011110000110101111111111101001100000100010100000000000100000111110101001101000001001111000001000001110100110100000111010100001100110100110011000100011101001101011111110111010000000000110100111111001100111101011111110001010011000111001101010101010011110000010001000111110001110111000000010001000111010101010001010000111101001101000100000111010011000100010111110011000001000101010011010011000000111101000100110001000100010011001100010101000111010111110100011111010011011101010111000000001111110001010000010111010100001101000001010000000100010000000001110001000100000000001101001111001100110001011101110011011101000101000011110000110111000011010001001101010101001101010100010111001101000101000000011101010111111100001101000011110000010011010101111111001101001100000000110111000000110001111111011101000101110001010100111100001101010011000000010000000100000000010100001111110000001100001101111100111100,2048'b11010011110011011101110100111100000101111100001100111111000001001111000101011111011111000001110101001100111101110111000100110000010111010101010100000101010011110100001101010101110011000100010011010000111100110101011101001111001100011101001101110111000011010001110101010000010000011101000101010101000111110111010001011111001111001101010101110001000000111100011101000100110100010101110001011111110001000011110100000001110100110000000011010011110100000000000101000101110101010111010111001101010000000100011101110111110100111101000011011111111100000011011100000000010001110000011101011100110000110000110111000100001101001101000000010001011100010101110001010011110000010100000100110101011101110000111100011101000001110111001101011100110001010001000100000011010001010011010000110000110111010011010011011100011100010100001101001100011101010111011100010000001101001101111100000101000111110011011100000100111100110011010100000000111101110111001100010000110000011100001101010011010000110001000000000000000011001100111100000000110100110011110011111111000101011101000000000011011100000101110100000011001101010100010000001100000000010100011100001111000100010100110000110101110011010101110100010101110100000011011111110100111111000001111111000011110101001111010011110101111111000100000000010001001111000011010100010100001111000011010111111100001100110001000100010100011101001101010101110111110000001101000101000111010111001100001101111100001100110011010111000101110100001101010101000001110101001100011101001101010011000101000001000100000101001111000101010000001101000000011100000001011111110001010001011111010001110100000000111101110000011101001111110101010000111100010100110011000000110101011101000111000001000111010011001100111111000100000001011100010011011100011100011111011111010001000100110011010000110101000000111111000000111100011111010100110111000011000100000111000011000011001100011100110100110001110000010101001111111100000001010101111100000000110111010000010100010011001101010100111111010000111100010101010000010000001100110011010000110000010111110111,2048'b00001111110001011100001111110011010011111101010011010011000100001101011111011111110111001101110111110100000111111101001100000011001111111101110000000111111111010011000001001100011101110000010101010001000001000001110100000101011101001111110011110101110011000000001111110001110101010000110101111100010011000000001111000001000011010101110001000100111111011100010011000001111101010100000100000101000000010101110001001100011101001100110100010001110111111111000001000100000000000000010011000000000000110100001101000111001111010101110000001100001111110101001101001111010111001101111111001111000101110011110000110111010111000101001111010100010001001100000001110001000001001111110001000100010111000100111101000101000001011111000111111101011111011100110000011101110001001100010100000001011100111111000101000000000111000001110001000001110011000000011100011111000100010111010111000111000101110100111111110111000100001111011100111100010000010001000001111111011101011101011101000101000001110111010100001111010011010011111101111111110000110000010001010101000111010111000101000000010011010000110011111101000111010101000111000111000001110100000100000000110100010111001101000001110100011101110011001100010100011111000111000011111111110011001111110100000101000011110100011111010001010000111111000101001100001111010111010001010100000100000011001101010111000100001100010011000000110001010101110100110000000000010100111111110011011100111101000101110000110000011111000100001100001101010001000000110111000100000000001111111101000100110101110011000111010000010011011101001100010100000000111111110111010011000011000111010100000001010100111100110001110001001101000001110111110111001101001100000011000100001100111100011100000101001100110001000101000100110101110000110111000001000111110101000100110001110000001101111111110100000011000000110001001100001111110001110000000100010000010001000011111111001100000101110011000000011101110000000000001111111111010100010001001100110011000011010101000101000101010100001100010000001100000111010100000101011101010101110101010000110001010000,2048'b01010001011100000101000111000100111111010100000001010011010101010000010100001100001111110100000001011100110111110101110011010001111100110011011100010101000111010100110000011100111111011100001111001101110011000000111100110111110001011100111101000111110101000100110000000001000000000100000001000101010011011101011101010111110101000001000011000000111111000100010000010000000111110000011100000111000100001111110011000100110011011101000101010100010011010100110101001100011100110100010000110001010001110101111101010100110000110011010101000111001111000101000100011111010111011111110011000111011101010100001101010100000000000111011100001111010100011101000001110001000100001100010100010111000001000000111100110101010101000100011111011101010111010011110000001101110011000000010111001101010101110111000001000111010111000001001100111101001100010100011101010111001111111100000000000011010100001100111100110001111100110111110101010101000100001101000100010101010001010100000000001101001100110100010100011111010000000111110100000011001111011111111100011100000001110101110000010000010100110000010111010001010000110101110100010100000111000000000101010011000101111100010111010011000011111101011101000000010001000011000001010001000111000101010000110011111111111100110100000001110001110100010000110100010001000101111101010011111111111111110011000100011101110011001101110000000000110000011100001111010111111101110111010000110101110001000011000000001100001100011111110111000011111111110101000101010000110001010011110111000001011100010111001101110001010111000011000001000000111101110011010001110011010000000100011100011101110101010111110100111101010000010100000011000101000000000100000000000000110000110000110100001111110101010000010000110000000001110000001100110011000000010001000100000011011100010000000001110101010111000101000011110000010000110000110100110111010111110000001100010000110011111101000111001101110100110000000111000011011101111100001101001101010111010100010100010000010100011100010101111100110101010111011111010100110011000111000101110011110101000000000100,2048'b11010011000000010100011100010011000101000001001111011101111100010100000100110001110100011101010011110100010011011101000001000100110001001101110100010000000011110000111111110100001101010011001100110100010000000000010101011111010111110000010001110100011101001111011111010000001100110111110000111100000001110111010011000100000100010001000000000001111111110011111101000011011101001100000000000101110100001100000011001111010101001100000100000111110011011100110111000000010000111111110100111100001100000011010001010000110101000011110011010101110001111100010001111100010011110101010001000100110000010101110001000111000111010101001101000111000100110000110100010000010011010111110001111111000011011111001101110000000100010100001100111111110011001111010000110101110000110001110111011101110100010111000001000000110011001100001100000101110111111101000111010101010011110100000100110100011100000001111111011101010001111101110000001101111111010101110000001111010000000111111100000001111101000011000000010000110001000111010011000100010000001111010111000111111100010101000011000111001100001100010100010001000100000001010011011100000000000011010100001111000000010001110001011101010101110011000100011101110101111100000001000001000111110011000100011101110100011101000111011100010000111101111111001101111111000000110011011111110101111111001101110100111111110111010101111100011100010111000101010000010000110101001101000001110101011101000011011101000111111100000100000011011100000101010100010001000100001101010011010101000111011101011111010011010101000111010111000100110101110000000100010001110100110000110000111100001101001100111100000111111101000011111100110001001100010100010011111101110101110000110000111100110011011111011101000001011100001100001100110000110000000000011100010101000111000100000111011101011111011101000101000111000100001100110011000000110111010111001100000011000001110100000011001101001111000000000011000001011101010100001111010100001100001101110000010100010100010001110011010011011111001100110011000101000101010000111100000101000000001101001100011101};
logic[127:0]weight_l3[9:0]={128'b01000101001111000011110001000100110001111101001100000101000000010000011100000000111100001101110101011111000100011111010111110001,128'b11111100110100111101010101000101110100010011000011110111110011111100111101010101110100110101111100010111010001111100110000111100,128'b11000011001100000001010001010011011111011101110100010100010100000001011111111111011100111111110001000011010001110011010011010100,128'b01010101110111010011001111110100110001000111010100010011000001001101010011110011001111011100000111001100110101001101010011000100,128'b00000000000101001101010100111111000111110001001101011100010111000011000000001111010001010011010101010001010001110000010011010101,128'b00000100000100000011001101010100010100000000001111000111000100000100010101110101000011110111011100001100001111010101010111011100,128'b00010011110000000000000000110011000111000100000011110100111101111111000101110000010111011111110000010111111101001100011111110000,128'b01000000111101011101001100000111110000011111010111111111000011001100110000011101110111110100010011111100010000000100000100000101,128'b01000111010101000001010000000001000100111101010001000000000000110011000011110011010000110011010000001101010000110111000001011101,128'b11000000110001010001111101110001010100010100000100010001011111110111010001011111110111110001110111000001111111010101000011110001};
logic[1:0]bias_l1[1023:0]={2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11};
logic[1:0]bias_l2[63:0]={2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11,2'b11};
logic[1:0]bias_l3[9:0]={2'b01,2'b01,2'b01,2'b01,2'b01,2'b01,2'b01,2'b01,2'b01,2'b01};
