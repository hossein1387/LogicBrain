../../CALCULATORUNIT/rtl/LineBufferL3.vhd