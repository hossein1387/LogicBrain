../../CALCULATORUNIT/rtl/AccelCoreL2.vhd