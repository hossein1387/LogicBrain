../../NEURALCORE/rtl/mega_ram.sv