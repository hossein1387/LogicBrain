../../CALCULATORUNIT/rtl/calculatorunit.sv