../../CALCULATORUNIT/rtl/AccelCoreL3.vhd