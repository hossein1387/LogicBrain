../../CALCULATORUNIT/rtl/PE.vhd